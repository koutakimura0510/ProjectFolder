
//
// Verific Verilog Description of module MTopTi180MIPI25GRxHDMIV101
//

module MTopTi180MIPI25GRxHDMIV101 (MipiDphyRx1_RESET_N, MipiDphyRx1_RST0_N, 
            MipiDphyRx1_STOPSTATE_CLK, MipiDphyRx1_STOPSTATE_LAN0, MipiDphyRx1_STOPSTATE_LAN1, 
            MipiDphyRx1_ERR_ESC_LAN0, MipiDphyRx1_ERR_ESC_LAN1, MipiDphyRx1_ERR_CONTROL_LAN0, 
            MipiDphyRx1_ERR_CONTROL_LAN1, MipiDphyRx1_TX_REQUEST_ESC, MipiDphyRx1_TURN_REQUEST, 
            MipiDphyRx1_FORCE_RX_MODE, MipiDphyRx1_TX_TRIGGER_ESC, MipiDphyRx1_RX_TRIGGER_ESC, 
            MipiDphyRx1_DIRECTION, MipiDphyRx1_ERR_CONTENTION_LP0, MipiDphyRx1_ERR_CONTENTION_LP1, 
            MipiDphyRx1_RX_CLK_ACTIVE_HS, MipiDphyRx1_RX_ACTIVE_HS_LAN0, 
            MipiDphyRx1_RX_ACTIVE_HS_LAN1, MipiDphyRx1_RX_VALID_HS_LAN0, 
            MipiDphyRx1_RX_VALID_HS_LAN1, MipiDphyRx1_RX_SYNC_HS_LAN0, MipiDphyRx1_RX_SYNC_HS_LAN1, 
            MipiDphyRx1_RX_SKEW_CAL_HS_LAN0, MipiDphyRx1_RX_SKEW_CAL_HS_LAN1, 
            MipiDphyRx1_RX_DATA_HS_LAN0, MipiDphyRx1_RX_DATA_HS_LAN1, MipiDphyRx1_ERR_SOT_HS_LAN0, 
            MipiDphyRx1_ERR_SOT_HS_LAN1, MipiDphyRx1_ERR_SOT_SYNC_HS_LAN0, 
            MipiDphyRx1_ERR_SOT_SYNC_HS_LAN1, MipiDphyRx1_RX_LPDT_ESC, MipiDphyRx1_RX_DATA_ESC, 
            MipiDphyRx1_RX_VALID_ESC, MipiDphyRx1_RX_ERR_SYNC_ESC, MipiDphyRx1_TX_LPDT_ESC, 
            MipiDphyRx1_TX_DATA_ESC, MipiDphyRx1_TX_VALID_ESC, MipiDphyRx1_TX_READY_ESC, 
            MipiDphyRx1_TX_ULPS_ESC, MipiDphyRx1_TX_ULPS_EXIT, MipiDphyRx1_RX_ULPS_CLK_NOT, 
            MipiDphyRx1_RX_ULPS_ACTIVE_CLK_NOT, MipiDphyRx1_RX_ULPS_ESC_LAN0, 
            MipiDphyRx1_RX_ULPS_ESC_LAN1, MipiDphyRx1_RX_ULPS_ACTIVE_NOT_LAN0, 
            MipiDphyRx1_RX_ULPS_ACTIVE_NOT_LAN1, MipiDphyRx1_WORD_CLKOUT_HS, 
            MipiDphyRx1_LP_CLK, MipiDphyRx1_RX_CLK_ESC_LAN0, MipiDphyRx1_RX_CLK_ESC_LAN1, 
            MipiDphyRx1_TX_CLK_ESC, oAdv7511Vs, oAdv7511Hs, oAdv7511De, 
            oAdv7511Data, iAdv7511Sda, oAdv7511SdaOe, iAdv7511Scl, oAdv7511SclOe, 
            oLed, iPushSw, iSCLK, iBCLK, iPCLK, iFCLK, pll_inst1_LOCKED, 
            pll_inst1_RSTN, iVCLK, pll_inst2_LOCKED, pll_inst2_RSTN, 
            pll_ddr_LOCKED, pll_ddr_RSTN, oTestPort, jtag_inst1_TDI, 
            jtag_inst1_TCK, jtag_inst1_TMS, jtag_inst1_TDO, jtag_inst1_SEL, 
            jtag_inst1_DRCK, jtag_inst1_RUNTEST, jtag_inst1_CAPTURE, jtag_inst1_SHIFT, 
            jtag_inst1_UPDATE, jtag_inst1_RESET, jtag_inst2_CAPTURE, jtag_inst2_DRCK, 
            jtag_inst2_RESET, jtag_inst2_RUNTEST, jtag_inst2_SEL, jtag_inst2_SHIFT, 
            jtag_inst2_TCK, jtag_inst2_TDI, jtag_inst2_TMS, jtag_inst2_UPDATE, 
            jtag_inst2_TDO);
    output MipiDphyRx1_RESET_N /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_RST0_N /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input MipiDphyRx1_STOPSTATE_CLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_STOPSTATE_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_STOPSTATE_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_ESC_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_ESC_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_CONTROL_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_CONTROL_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output MipiDphyRx1_TX_REQUEST_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_TURN_REQUEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_FORCE_RX_MODE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [3:0]MipiDphyRx1_TX_TRIGGER_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input [3:0]MipiDphyRx1_RX_TRIGGER_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_DIRECTION /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_CONTENTION_LP0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_CONTENTION_LP1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_CLK_ACTIVE_HS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ACTIVE_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ACTIVE_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_VALID_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_VALID_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_SYNC_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_SYNC_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_SKEW_CAL_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_SKEW_CAL_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]MipiDphyRx1_RX_DATA_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]MipiDphyRx1_RX_DATA_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_SOT_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_SOT_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_SOT_SYNC_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_SOT_SYNC_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_LPDT_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]MipiDphyRx1_RX_DATA_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_VALID_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ERR_SYNC_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output MipiDphyRx1_TX_LPDT_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]MipiDphyRx1_TX_DATA_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_TX_VALID_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_TX_READY_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_TX_ULPS_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_TX_ULPS_EXIT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_CLK_NOT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ACTIVE_CLK_NOT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ESC_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ESC_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ACTIVE_NOT_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ACTIVE_NOT_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_WORD_CLKOUT_HS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_LP_CLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_CLK_ESC_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_CLK_ESC_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output MipiDphyRx1_TX_CLK_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output oAdv7511Vs /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output oAdv7511Hs /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output oAdv7511De /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [15:0]oAdv7511Data /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input iAdv7511Sda /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output oAdv7511SdaOe /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input iAdv7511Scl /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output oAdv7511SclOe /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [5:0]oLed /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input [1:0]iPushSw /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input iSCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input iBCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input iPCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input iFCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input pll_inst1_LOCKED /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output pll_inst1_RSTN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input iVCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input pll_inst2_LOCKED /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output pll_inst2_RSTN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input pll_ddr_LOCKED /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output pll_ddr_RSTN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [25:0]oTestPort /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input jtag_inst1_TDI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TMS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output jtag_inst1_TDO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input jtag_inst1_SEL /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_DRCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RUNTEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_CAPTURE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SHIFT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_UPDATE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RESET /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_CAPTURE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_DRCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_RESET /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_RUNTEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_SEL /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_SHIFT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_TCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_TDI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_TMS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_UPDATE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output jtag_inst2_TDO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    
    wire la0_probe4, la0_probe10, rFRST, rBRST, rVRST, rnVRST, la0_probe2, 
        la0_probe11, \la0_probe6[0] , \la0_probe9[0] , \MCsiRxController/MCsi2Decoder/rHsSt[0] , 
        \la0_probe3[0] , \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd , 
        la0_probe5, la0_probe7, n117, n118, la0_probe0, n120, n121, 
        \MCsiRxController/wHsPixel[0] , \MCsiRxController/MCsi2Decoder/wFtiRvd[0] , 
        n124, n125, \MCsiRxController/wHsValid , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] , 
        \MCsiRxController/MCsi2Decoder/rHsSt[2] , \MCsiRxController/MCsi2Decoder/rHsSt[1] , 
        \la0_probe9[7] , \la0_probe9[6] , \la0_probe9[5] , \la0_probe9[4] , 
        \la0_probe9[3] , \la0_probe9[2] , \la0_probe9[1] , \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] , 
        \MCsiRxController/MCsi2Decoder/wFtiEmp[0] , \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] , 
        n169, n170, \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[16] , n189, n190, \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9] , 
        n210, n211, \MCsiRxController/wHsPixel[1] , \MCsiRxController/wHsPixel[2] , 
        \MCsiRxController/wHsPixel[3] , \MCsiRxController/wHsPixel[4] , 
        \MCsiRxController/wHsPixel[5] , \MCsiRxController/wHsPixel[6] , 
        \MCsiRxController/wHsPixel[7] , \MCsiRxController/wHsPixel[8] , 
        \MCsiRxController/wHsPixel[9] , \MCsiRxController/wHsPixel[10] , 
        \MCsiRxController/wHsPixel[11] , \MCsiRxController/wHsPixel[12] , 
        \MCsiRxController/wHsPixel[13] , \MCsiRxController/wHsPixel[14] , 
        \MCsiRxController/wHsPixel[15] , \wHsWordCnt[1] , \wHsWordCnt[2] , 
        \wHsWordCnt[3] , \wHsWordCnt[4] , \wHsWordCnt[5] , \wHsWordCnt[6] , 
        \wHsWordCnt[7] , \wHsWordCnt[8] , \wHsWordCnt[9] , \wHsWordCnt[10] , 
        \wHsWordCnt[11] , \wHsWordCnt[12] , \wHsWordCnt[13] , \wHsWordCnt[14] , 
        \wHsWordCnt[15] , \wHsDatatype[2] , \wHsDatatype[3] , \wHsDatatype[4] , 
        \wHsDatatype[5] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12] , \la0_probe8[0] , 
        \la0_probe8[1] , \la0_probe8[2] , \la0_probe8[3] , \la0_probe8[4] , 
        \la0_probe8[5] , \la0_probe8[6] , \la0_probe8[7] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0] , wVideoVd, n295, 
        n296, \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] , \MCsiRxController/wFtiEmp[0] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1] , \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3] , \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5] , \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7] , \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8] , 
        \wVideoPixel[0] , \wVideoPixel[1] , \wVideoPixel[2] , \wVideoPixel[3] , 
        \wVideoPixel[4] , \wVideoPixel[5] , \wVideoPixel[6] , \wVideoPixel[7] , 
        \wVideoPixel[8] , \wVideoPixel[9] , \wVideoPixel[10] , \wVideoPixel[11] , 
        \wVideoPixel[12] , \wVideoPixel[13] , \wVideoPixel[14] , \wVideoPixel[15] , 
        n331, n332, \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] , 
        \la0_probe6[1] , \la0_probe6[2] , \la0_probe6[3] , \la0_probe6[4] , 
        \la0_probe6[5] , \la0_probe6[6] , \la0_probe6[7] , \la0_probe6[8] , 
        \la0_probe6[9] , \la0_probe6[10] , \la0_probe6[11] , \la0_probe6[12] , 
        \la0_probe6[13] , \la0_probe6[14] , \la0_probe6[15] , \la0_probe3[1] , 
        \MVideoPostProcess/rVtgRstCnt[0] , \MVideoPostProcess/rVtgRST[0] , 
        \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] , \MVideoPostProcess/inst_adv7511_config/r_m_en_1P , 
        \MVideoPostProcess/inst_adv7511_config/r_last_1P , \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] , \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0] , \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P , \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] , 
        \MVideoPostProcess/inst_adv7511_config/w_ack , \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] , 
        \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[0] , n436, n437, 
        \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[1] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[2] , 
        \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[3] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[4] , 
        \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[5] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[6] , 
        \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[7] , \MVideoPostProcess/mVideoTimingGen/dff_27/i4_pre , 
        \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0 , \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3 , 
        \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] , 
        \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] , 
        \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] , 
        \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14] , 
        \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] , \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3] , \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] , 
        \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] , \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6] , 
        \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7] , \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1] , 
        \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2] , \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3] , 
        \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4] , \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5] , 
        \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6] , \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7] , 
        \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] , 
        n492, n493, \MVideoPostProcess/mVideoTimingGen/rVpos[0] , n495, 
        n496, \MVideoPostProcess/mVideoTimingGen/rVde[0] , \MVideoPostProcess/mVideoTimingGen/rHpos[0] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[1] , \MVideoPostProcess/mVideoTimingGen/rVpos[2] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[3] , \MVideoPostProcess/mVideoTimingGen/rVpos[4] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[5] , \MVideoPostProcess/mVideoTimingGen/rVpos[6] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[7] , \MVideoPostProcess/mVideoTimingGen/rVpos[8] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[9] , \MVideoPostProcess/mVideoTimingGen/rVpos[10] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[11] , \MVideoPostProcess/mVideoTimingGen/dff_11/i4_pre , 
        \MVideoPostProcess/mVideoTimingGen/rVde[1] , \MVideoPostProcess/mVideoTimingGen/rVde[3] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[1] , \MVideoPostProcess/mVideoTimingGen/rHpos[2] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[3] , \MVideoPostProcess/mVideoTimingGen/rHpos[4] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[5] , \MVideoPostProcess/mVideoTimingGen/rHpos[6] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[7] , \MVideoPostProcess/mVideoTimingGen/rHpos[8] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[9] , \MVideoPostProcess/mVideoTimingGen/rHpos[10] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0] , 
        wVideofull, n532, n533, \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12] , 
        n560, n561, \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0] , 
        n577, n578, \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12] , 
        n604, n605, \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0] , 
        n621, n622, \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12] , 
        n648, n649, \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0] , 
        n665, n666, \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12] , 
        n692, n693, \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0] , 
        n709, n710, \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12] , 
        n736, n737, \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0] , 
        n753, n754, \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12] , 
        n780, n781, \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0] , 
        n797, n798, \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12] , 
        n824, n825, \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0] , 
        n841, n842, \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12] , 
        n868, n869, \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0] , 
        n885, n886, \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12] , 
        n912, n913, \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0] , 
        n929, n930, \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12] , 
        n956, n957, \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0] , 
        n973, n974, \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12] , 
        n1000, n1001, \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0] , 
        n1017, n1018, \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12] , 
        n1044, n1045, \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0] , 
        n1061, n1062, \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12] , 
        n1088, n1089, \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0] , 
        n1105, n1106, \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12] , 
        n1132, n1133, \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0] , 
        n1149, n1150, \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12] , 
        n1176, n1177, \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0] , 
        n1193, \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12] , 
        n1219, n1220, \MVideoPostProcess/rVtgRstCnt[1] , \MVideoPostProcess/rVtgRstCnt[2] , 
        \MVideoPostProcess/rVtgRstCnt[3] , \MVideoPostProcess/rVtgRstCnt[4] , 
        \MVideoPostProcess/rVtgRstCnt[5] , \MVideoPostProcess/rVtgRstCnt[6] , 
        \MVideoPostProcess/rVtgRstCnt[7] , \MVideoPostProcess/rVtgRstCnt[8] , 
        \MVideoPostProcess/rVtgRstCnt[9] , \MVideoPostProcess/rVtgRstCnt[10] , 
        \MVideoPostProcess/rVtgRST[1] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] , 
        \genblk1.genblk1[0].mPulseGenerator/rSft[0] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[12] , \genblk1.genblk1[0].mPulseGenerator/rSft[1] , 
        \genblk1.genblk1[0].mPulseGenerator/rSft[2] , \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0] , 
        \genblk1.genblk1[3].mPulseGenerator/rSft[0] , \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] , 
        \genblk1.genblk1[3].mPulseGenerator/rSft[1] , \genblk1.genblk1[3].mPulseGenerator/rSft[2] , 
        \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0] , \genblk1.genblk1[4].mPulseGenerator/rSft[0] , 
        \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] , \genblk1.genblk1[4].mPulseGenerator/rSft[1] , 
        \genblk1.genblk1[4].mPulseGenerator/rSft[2] , \edb_top_inst/n2759 , 
        \edb_top_inst/la0/la_run_trig , \edb_top_inst/la0/la_trig_pattern[0] , 
        \edb_top_inst/la0/la_run_trig_imdt , \edb_top_inst/la0/la_stop_trig , 
        \edb_top_inst/la0/la_capture_pattern[0] , \edb_top_inst/la0/la_trig_mask[0] , 
        \edb_top_inst/la0/la_num_trigger[0] , \edb_top_inst/la0/la_window_depth[0] , 
        \edb_top_inst/la0/la_soft_reset_in , \edb_top_inst/la0/address_counter[0] , 
        \edb_top_inst/la0/opcode[0] , \edb_top_inst/la0/bit_count[0] , \edb_top_inst/la0/word_count[0] , 
        \edb_top_inst/la0/data_out_shift_reg[0] , \edb_top_inst/la0/module_state[0] , 
        \edb_top_inst/la0/la_resetn_p1 , \edb_top_inst/la0/la_resetn , \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/cap_fifo_din_cu[0] , \edb_top_inst/la0/cap_fifo_din_tu[0] , 
        \edb_top_inst/la0/internal_register_select[0] , \edb_top_inst/la0/la_trig_pos[0] , 
        \edb_top_inst/la0/la_trig_pattern[1] , \edb_top_inst/la0/la_capture_pattern[1] , 
        \edb_top_inst/la0/la_trig_mask[1] , \edb_top_inst/la0/la_trig_mask[2] , 
        \edb_top_inst/la0/la_trig_mask[3] , \edb_top_inst/la0/la_trig_mask[4] , 
        \edb_top_inst/la0/la_trig_mask[5] , \edb_top_inst/la0/la_trig_mask[6] , 
        \edb_top_inst/la0/la_trig_mask[7] , \edb_top_inst/la0/la_trig_mask[8] , 
        \edb_top_inst/la0/la_trig_mask[9] , \edb_top_inst/la0/la_trig_mask[10] , 
        \edb_top_inst/la0/la_trig_mask[11] , \edb_top_inst/la0/la_trig_mask[12] , 
        \edb_top_inst/la0/la_trig_mask[13] , \edb_top_inst/la0/la_trig_mask[14] , 
        \edb_top_inst/la0/la_trig_mask[15] , \edb_top_inst/la0/la_trig_mask[16] , 
        \edb_top_inst/la0/la_trig_mask[17] , \edb_top_inst/la0/la_trig_mask[18] , 
        \edb_top_inst/la0/la_trig_mask[19] , \edb_top_inst/la0/la_trig_mask[20] , 
        \edb_top_inst/la0/la_trig_mask[21] , \edb_top_inst/la0/la_trig_mask[22] , 
        \edb_top_inst/la0/la_trig_mask[23] , \edb_top_inst/la0/la_trig_mask[24] , 
        \edb_top_inst/la0/la_trig_mask[25] , \edb_top_inst/la0/la_trig_mask[26] , 
        \edb_top_inst/la0/la_trig_mask[27] , \edb_top_inst/la0/la_trig_mask[28] , 
        \edb_top_inst/la0/la_trig_mask[29] , \edb_top_inst/la0/la_trig_mask[30] , 
        \edb_top_inst/la0/la_trig_mask[31] , \edb_top_inst/la0/la_trig_mask[32] , 
        \edb_top_inst/la0/la_trig_mask[33] , \edb_top_inst/la0/la_trig_mask[34] , 
        \edb_top_inst/la0/la_trig_mask[35] , \edb_top_inst/la0/la_trig_mask[36] , 
        \edb_top_inst/la0/la_trig_mask[37] , \edb_top_inst/la0/la_trig_mask[38] , 
        \edb_top_inst/la0/la_trig_mask[39] , \edb_top_inst/la0/la_trig_mask[40] , 
        \edb_top_inst/la0/la_trig_mask[41] , \edb_top_inst/la0/la_trig_mask[42] , 
        \edb_top_inst/la0/la_trig_mask[43] , \edb_top_inst/la0/la_trig_mask[44] , 
        \edb_top_inst/la0/la_trig_mask[45] , \edb_top_inst/la0/la_trig_mask[46] , 
        \edb_top_inst/la0/la_trig_mask[47] , \edb_top_inst/la0/la_trig_mask[48] , 
        \edb_top_inst/la0/la_trig_mask[49] , \edb_top_inst/la0/la_trig_mask[50] , 
        \edb_top_inst/la0/la_trig_mask[51] , \edb_top_inst/la0/la_trig_mask[52] , 
        \edb_top_inst/la0/la_trig_mask[53] , \edb_top_inst/la0/la_trig_mask[54] , 
        \edb_top_inst/la0/la_trig_mask[55] , \edb_top_inst/la0/la_trig_mask[56] , 
        \edb_top_inst/la0/la_trig_mask[57] , \edb_top_inst/la0/la_trig_mask[58] , 
        \edb_top_inst/la0/la_trig_mask[59] , \edb_top_inst/la0/la_trig_mask[60] , 
        \edb_top_inst/la0/la_trig_mask[61] , \edb_top_inst/la0/la_trig_mask[62] , 
        \edb_top_inst/la0/la_trig_mask[63] , \edb_top_inst/la0/la_num_trigger[1] , 
        \edb_top_inst/la0/la_num_trigger[2] , \edb_top_inst/la0/la_num_trigger[3] , 
        \edb_top_inst/la0/la_num_trigger[4] , \edb_top_inst/la0/la_num_trigger[5] , 
        \edb_top_inst/la0/la_num_trigger[6] , \edb_top_inst/la0/la_num_trigger[7] , 
        \edb_top_inst/la0/la_num_trigger[8] , \edb_top_inst/la0/la_num_trigger[9] , 
        \edb_top_inst/la0/la_num_trigger[10] , \edb_top_inst/la0/la_num_trigger[11] , 
        \edb_top_inst/la0/la_num_trigger[12] , \edb_top_inst/la0/la_num_trigger[13] , 
        \edb_top_inst/la0/la_num_trigger[14] , \edb_top_inst/la0/la_num_trigger[15] , 
        \edb_top_inst/la0/la_num_trigger[16] , \edb_top_inst/la0/la_window_depth[1] , 
        \edb_top_inst/la0/la_window_depth[2] , \edb_top_inst/la0/la_window_depth[3] , 
        \edb_top_inst/la0/la_window_depth[4] , \edb_top_inst/la0/address_counter[1] , 
        \edb_top_inst/la0/address_counter[2] , \edb_top_inst/la0/address_counter[3] , 
        \edb_top_inst/la0/address_counter[4] , \edb_top_inst/la0/address_counter[5] , 
        \edb_top_inst/la0/address_counter[6] , \edb_top_inst/la0/address_counter[7] , 
        \edb_top_inst/la0/address_counter[8] , \edb_top_inst/la0/address_counter[9] , 
        \edb_top_inst/la0/address_counter[10] , \edb_top_inst/la0/address_counter[11] , 
        \edb_top_inst/la0/address_counter[12] , \edb_top_inst/la0/address_counter[13] , 
        \edb_top_inst/la0/address_counter[14] , \edb_top_inst/la0/address_counter[15] , 
        \edb_top_inst/la0/address_counter[16] , \edb_top_inst/la0/address_counter[17] , 
        \edb_top_inst/la0/address_counter[18] , \edb_top_inst/la0/address_counter[19] , 
        \edb_top_inst/la0/address_counter[20] , \edb_top_inst/la0/address_counter[21] , 
        \edb_top_inst/la0/address_counter[22] , \edb_top_inst/la0/address_counter[23] , 
        \edb_top_inst/la0/address_counter[24] , \edb_top_inst/la0/address_counter[25] , 
        \edb_top_inst/la0/address_counter[26] , \edb_top_inst/la0/opcode[1] , 
        \edb_top_inst/la0/opcode[2] , \edb_top_inst/la0/opcode[3] , \edb_top_inst/la0/bit_count[1] , 
        \edb_top_inst/la0/bit_count[2] , \edb_top_inst/la0/bit_count[3] , 
        \edb_top_inst/la0/bit_count[4] , \edb_top_inst/la0/bit_count[5] , 
        \edb_top_inst/la0/word_count[1] , \edb_top_inst/la0/word_count[2] , 
        \edb_top_inst/la0/word_count[3] , \edb_top_inst/la0/word_count[4] , 
        \edb_top_inst/la0/word_count[5] , \edb_top_inst/la0/word_count[6] , 
        \edb_top_inst/la0/word_count[7] , \edb_top_inst/la0/word_count[8] , 
        \edb_top_inst/la0/word_count[9] , \edb_top_inst/la0/word_count[10] , 
        \edb_top_inst/la0/word_count[11] , \edb_top_inst/la0/word_count[12] , 
        \edb_top_inst/la0/word_count[13] , \edb_top_inst/la0/word_count[14] , 
        \edb_top_inst/la0/word_count[15] , \edb_top_inst/la0/data_out_shift_reg[1] , 
        \edb_top_inst/la0/data_out_shift_reg[2] , \edb_top_inst/la0/data_out_shift_reg[3] , 
        \edb_top_inst/la0/data_out_shift_reg[4] , \edb_top_inst/la0/data_out_shift_reg[5] , 
        \edb_top_inst/la0/data_out_shift_reg[6] , \edb_top_inst/la0/data_out_shift_reg[7] , 
        \edb_top_inst/la0/data_out_shift_reg[8] , \edb_top_inst/la0/data_out_shift_reg[9] , 
        \edb_top_inst/la0/data_out_shift_reg[10] , \edb_top_inst/la0/data_out_shift_reg[11] , 
        \edb_top_inst/la0/data_out_shift_reg[12] , \edb_top_inst/la0/data_out_shift_reg[13] , 
        \edb_top_inst/la0/data_out_shift_reg[14] , \edb_top_inst/la0/data_out_shift_reg[15] , 
        \edb_top_inst/la0/data_out_shift_reg[16] , \edb_top_inst/la0/data_out_shift_reg[17] , 
        \edb_top_inst/la0/data_out_shift_reg[18] , \edb_top_inst/la0/data_out_shift_reg[19] , 
        \edb_top_inst/la0/data_out_shift_reg[20] , \edb_top_inst/la0/data_out_shift_reg[21] , 
        \edb_top_inst/la0/data_out_shift_reg[22] , \edb_top_inst/la0/data_out_shift_reg[23] , 
        \edb_top_inst/la0/data_out_shift_reg[24] , \edb_top_inst/la0/data_out_shift_reg[25] , 
        \edb_top_inst/la0/data_out_shift_reg[26] , \edb_top_inst/la0/data_out_shift_reg[27] , 
        \edb_top_inst/la0/data_out_shift_reg[28] , \edb_top_inst/la0/data_out_shift_reg[29] , 
        \edb_top_inst/la0/data_out_shift_reg[30] , \edb_top_inst/la0/data_out_shift_reg[31] , 
        \edb_top_inst/la0/data_out_shift_reg[32] , \edb_top_inst/la0/data_out_shift_reg[33] , 
        \edb_top_inst/la0/data_out_shift_reg[34] , \edb_top_inst/la0/data_out_shift_reg[35] , 
        \edb_top_inst/la0/data_out_shift_reg[36] , \edb_top_inst/la0/data_out_shift_reg[37] , 
        \edb_top_inst/la0/data_out_shift_reg[38] , \edb_top_inst/la0/data_out_shift_reg[39] , 
        \edb_top_inst/la0/data_out_shift_reg[40] , \edb_top_inst/la0/data_out_shift_reg[41] , 
        \edb_top_inst/la0/data_out_shift_reg[42] , \edb_top_inst/la0/data_out_shift_reg[43] , 
        \edb_top_inst/la0/data_out_shift_reg[44] , \edb_top_inst/la0/data_out_shift_reg[45] , 
        \edb_top_inst/la0/data_out_shift_reg[46] , \edb_top_inst/la0/data_out_shift_reg[47] , 
        \edb_top_inst/la0/data_out_shift_reg[48] , \edb_top_inst/la0/data_out_shift_reg[49] , 
        \edb_top_inst/la0/data_out_shift_reg[50] , \edb_top_inst/la0/data_out_shift_reg[51] , 
        \edb_top_inst/la0/data_out_shift_reg[52] , \edb_top_inst/la0/data_out_shift_reg[53] , 
        \edb_top_inst/la0/data_out_shift_reg[54] , \edb_top_inst/la0/data_out_shift_reg[55] , 
        \edb_top_inst/la0/data_out_shift_reg[56] , \edb_top_inst/la0/data_out_shift_reg[57] , 
        \edb_top_inst/la0/data_out_shift_reg[58] , \edb_top_inst/la0/data_out_shift_reg[59] , 
        \edb_top_inst/la0/data_out_shift_reg[60] , \edb_top_inst/la0/data_out_shift_reg[61] , 
        \edb_top_inst/la0/data_out_shift_reg[62] , \edb_top_inst/la0/data_out_shift_reg[63] , 
        \edb_top_inst/la0/module_state[1] , \edb_top_inst/la0/module_state[2] , 
        \edb_top_inst/la0/module_state[3] , \edb_top_inst/la0/crc_data_out[0] , 
        \edb_top_inst/la0/crc_data_out[1] , \edb_top_inst/la0/crc_data_out[2] , 
        \edb_top_inst/la0/crc_data_out[3] , \edb_top_inst/la0/crc_data_out[4] , 
        \edb_top_inst/la0/crc_data_out[5] , \edb_top_inst/la0/crc_data_out[6] , 
        \edb_top_inst/la0/crc_data_out[7] , \edb_top_inst/la0/crc_data_out[8] , 
        \edb_top_inst/la0/crc_data_out[9] , \edb_top_inst/la0/crc_data_out[10] , 
        \edb_top_inst/la0/crc_data_out[11] , \edb_top_inst/la0/crc_data_out[12] , 
        \edb_top_inst/la0/crc_data_out[13] , \edb_top_inst/la0/crc_data_out[14] , 
        \edb_top_inst/la0/crc_data_out[15] , \edb_top_inst/la0/crc_data_out[16] , 
        \edb_top_inst/la0/crc_data_out[17] , \edb_top_inst/la0/crc_data_out[18] , 
        \edb_top_inst/la0/crc_data_out[19] , \edb_top_inst/la0/crc_data_out[20] , 
        \edb_top_inst/la0/crc_data_out[21] , \edb_top_inst/la0/crc_data_out[22] , 
        \edb_top_inst/la0/crc_data_out[23] , \edb_top_inst/la0/crc_data_out[24] , 
        \edb_top_inst/la0/crc_data_out[25] , \edb_top_inst/la0/crc_data_out[26] , 
        \edb_top_inst/la0/crc_data_out[27] , \edb_top_inst/la0/crc_data_out[28] , 
        \edb_top_inst/la0/crc_data_out[29] , \edb_top_inst/la0/crc_data_out[30] , 
        \edb_top_inst/la0/crc_data_out[31] , \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout , \edb_top_inst/la0/tu_trigger , 
        \edb_top_inst/la0/cap_fifo_din_cu[1] , \edb_top_inst/la0/cap_fifo_din_cu[2] , 
        \edb_top_inst/la0/cap_fifo_din_cu[5] , \edb_top_inst/la0/cap_fifo_din_cu[6] , 
        \edb_top_inst/la0/cap_fifo_din_cu[23] , \edb_top_inst/la0/cap_fifo_din_cu[40] , 
        \edb_top_inst/la0/cap_fifo_din_cu[41] , \edb_top_inst/la0/cap_fifo_din_tu[1] , 
        \edb_top_inst/la0/cap_fifo_din_tu[2] , \edb_top_inst/la0/cap_fifo_din_tu[5] , 
        \edb_top_inst/la0/cap_fifo_din_tu[6] , \edb_top_inst/la0/cap_fifo_din_tu[23] , 
        \edb_top_inst/la0/cap_fifo_din_tu[40] , \edb_top_inst/la0/cap_fifo_din_tu[41] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[0] , \edb_top_inst/la0/la_biu_inst/run_trig_p2 , 
        \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 , \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 , 
        \edb_top_inst/la0/la_biu_inst/str_sync , \edb_top_inst/la0/la_biu_inst/str_sync_wbff1 , 
        \edb_top_inst/la0/la_biu_inst/str_sync_wbff2 , \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync , \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 , \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q , 
        \edb_top_inst/la0/data_from_biu[0] , \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[3] , \edb_top_inst/la0/la_biu_inst/curr_state[2] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[1] , \edb_top_inst/la0/biu_ready , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[15] , \edb_top_inst/la0/la_biu_inst/addr_reg[16] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[17] , \edb_top_inst/la0/la_biu_inst/addr_reg[18] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[19] , \edb_top_inst/la0/la_biu_inst/addr_reg[20] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[21] , \edb_top_inst/la0/la_biu_inst/addr_reg[22] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[23] , \edb_top_inst/la0/la_biu_inst/addr_reg[24] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[25] , \edb_top_inst/la0/la_biu_inst/addr_reg[26] , 
        \edb_top_inst/la0/data_from_biu[1] , \edb_top_inst/la0/data_from_biu[2] , 
        \edb_top_inst/la0/data_from_biu[3] , \edb_top_inst/la0/data_from_biu[4] , 
        \edb_top_inst/la0/data_from_biu[5] , \edb_top_inst/la0/data_from_biu[6] , 
        \edb_top_inst/la0/data_from_biu[7] , \edb_top_inst/la0/data_from_biu[8] , 
        \edb_top_inst/la0/data_from_biu[9] , \edb_top_inst/la0/data_from_biu[10] , 
        \edb_top_inst/la0/data_from_biu[11] , \edb_top_inst/la0/data_from_biu[12] , 
        \edb_top_inst/la0/data_from_biu[13] , \edb_top_inst/la0/data_from_biu[14] , 
        \edb_top_inst/la0/data_from_biu[15] , \edb_top_inst/la0/data_from_biu[16] , 
        \edb_top_inst/la0/data_from_biu[17] , \edb_top_inst/la0/data_from_biu[18] , 
        \edb_top_inst/la0/data_from_biu[19] , \edb_top_inst/la0/data_from_biu[20] , 
        \edb_top_inst/la0/data_from_biu[21] , \edb_top_inst/la0/data_from_biu[22] , 
        \edb_top_inst/la0/data_from_biu[23] , \edb_top_inst/la0/data_from_biu[24] , 
        \edb_top_inst/la0/data_from_biu[25] , \edb_top_inst/la0/data_from_biu[26] , 
        \edb_top_inst/la0/data_from_biu[27] , \edb_top_inst/la0/data_from_biu[28] , 
        \edb_top_inst/la0/data_from_biu[29] , \edb_top_inst/la0/data_from_biu[30] , 
        \edb_top_inst/la0/data_from_biu[31] , \edb_top_inst/la0/data_from_biu[32] , 
        \edb_top_inst/la0/data_from_biu[33] , \edb_top_inst/la0/data_from_biu[34] , 
        \edb_top_inst/la0/data_from_biu[35] , \edb_top_inst/la0/data_from_biu[36] , 
        \edb_top_inst/la0/data_from_biu[37] , \edb_top_inst/la0/data_from_biu[38] , 
        \edb_top_inst/la0/data_from_biu[39] , \edb_top_inst/la0/data_from_biu[40] , 
        \edb_top_inst/la0/data_from_biu[41] , \edb_top_inst/la0/data_from_biu[42] , 
        \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] , 
        \edb_top_inst/la0/la_sample_cnt[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[0] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] , 
        \edb_top_inst/la0/la_sample_cnt[1] , \edb_top_inst/la0/la_sample_cnt[2] , 
        \edb_top_inst/la0/la_sample_cnt[3] , \edb_top_inst/la0/la_sample_cnt[4] , 
        \edb_top_inst/la0/la_sample_cnt[5] , \edb_top_inst/la0/la_sample_cnt[6] , 
        \edb_top_inst/la0/la_sample_cnt[7] , \edb_top_inst/la0/la_sample_cnt[8] , 
        \edb_top_inst/la0/la_sample_cnt[9] , \edb_top_inst/la0/la_sample_cnt[10] , 
        \edb_top_inst/la0/la_sample_cnt[11] , \edb_top_inst/la0/la_sample_cnt[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[1] , \edb_top_inst/la0/la_biu_inst/fifo_counter[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[3] , \edb_top_inst/la0/la_biu_inst/fifo_counter[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[5] , \edb_top_inst/la0/la_biu_inst/fifo_counter[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[7] , \edb_top_inst/la0/la_biu_inst/fifo_counter[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[9] , \edb_top_inst/la0/la_biu_inst/fifo_counter[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[11] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] , 
        \edb_top_inst/la0/internal_register_select[1] , \edb_top_inst/la0/internal_register_select[2] , 
        \edb_top_inst/la0/internal_register_select[3] , \edb_top_inst/la0/internal_register_select[4] , 
        \edb_top_inst/la0/internal_register_select[5] , \edb_top_inst/la0/internal_register_select[6] , 
        \edb_top_inst/la0/internal_register_select[7] , \edb_top_inst/la0/internal_register_select[8] , 
        \edb_top_inst/la0/internal_register_select[9] , \edb_top_inst/la0/internal_register_select[10] , 
        \edb_top_inst/la0/internal_register_select[11] , \edb_top_inst/la0/internal_register_select[12] , 
        \edb_top_inst/la0/la_trig_pos[1] , \edb_top_inst/la0/la_trig_pos[2] , 
        \edb_top_inst/la0/la_trig_pos[3] , \edb_top_inst/la0/la_trig_pos[4] , 
        \edb_top_inst/la0/la_trig_pos[5] , \edb_top_inst/la0/la_trig_pos[6] , 
        \edb_top_inst/la0/la_trig_pos[7] , \edb_top_inst/la0/la_trig_pos[8] , 
        \edb_top_inst/la0/la_trig_pos[9] , \edb_top_inst/la0/la_trig_pos[10] , 
        \edb_top_inst/la0/la_trig_pos[11] , \edb_top_inst/la0/la_trig_pos[12] , 
        \edb_top_inst/la0/la_trig_pos[13] , \edb_top_inst/la0/la_trig_pos[14] , 
        \edb_top_inst/la0/la_trig_pos[15] , \edb_top_inst/la0/la_trig_pos[16] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[0] , \edb_top_inst/debug_hub_inst/module_id_reg[1] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[2] , \edb_top_inst/debug_hub_inst/module_id_reg[3] , 
        \edb_top_inst/n68 , \edb_top_inst/n70 , \edb_top_inst/n74 , \edb_top_inst/n694 , 
        \edb_top_inst/n696 , \edb_top_inst/n697 , \edb_top_inst/n698 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i40_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i35_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i36_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i37_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i38_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i39_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_pre , 
        \edb_top_inst/n2760 , \edb_top_inst/n2761 , \edb_top_inst/n2762 , 
        \edb_top_inst/n2763 , \edb_top_inst/n2764 , \edb_top_inst/n2765 , 
        \edb_top_inst/n2766 , \edb_top_inst/n2767 , \edb_top_inst/n2768 , 
        \edb_top_inst/n2769 , \edb_top_inst/n2770 , \edb_top_inst/n2771 , 
        \edb_top_inst/n2772 , \edb_top_inst/n2773 , \edb_top_inst/n2774 , 
        \edb_top_inst/n2775 , \edb_top_inst/n2776 , \edb_top_inst/n2777 , 
        \edb_top_inst/n2778 , \edb_top_inst/n2779 , \edb_top_inst/n2780 , 
        \edb_top_inst/n2781 , \edb_top_inst/n2782 , \edb_top_inst/n2783 , 
        \edb_top_inst/n2784 , \edb_top_inst/n2785 , \edb_top_inst/n2786 , 
        \edb_top_inst/n2787 , \edb_top_inst/n2788 , \edb_top_inst/n2789 , 
        \edb_top_inst/n2790 , \edb_top_inst/n2791 , \edb_top_inst/n2792 , 
        \edb_top_inst/n2793 , \edb_top_inst/n2794 , \edb_top_inst/n2795 , 
        \edb_top_inst/n2796 , \edb_top_inst/n2797 , \edb_top_inst/n2798 , 
        \edb_top_inst/n2799 , \edb_top_inst/n2800 , \edb_top_inst/n2801 , 
        \edb_top_inst/n2802 , \edb_top_inst/n2803 , \edb_top_inst/n2804 , 
        \edb_top_inst/n2805 , \edb_top_inst/n2806 , \edb_top_inst/n2807 , 
        \edb_top_inst/n2808 , \edb_top_inst/n2809 , \edb_top_inst/n2810 , 
        \edb_top_inst/n2811 , \edb_top_inst/n2812 , \edb_top_inst/n2813 , 
        \edb_top_inst/n2814 , \edb_top_inst/n2815 , \edb_top_inst/n2816 , 
        \edb_top_inst/n2817 , \edb_top_inst/n2818 , \edb_top_inst/n2819 , 
        \edb_top_inst/n2820 , \edb_top_inst/n2736 , \edb_top_inst/n2733 , 
        \edb_top_inst/n2821 , \edb_top_inst/n1249 , \edb_top_inst/n2822 , 
        \edb_top_inst/n2823 , \edb_top_inst/n2824 , \edb_top_inst/n2825 , 
        \edb_top_inst/n2826 , \edb_top_inst/n2827 , \edb_top_inst/n2828 , 
        \edb_top_inst/n2829 , \edb_top_inst/n2830 , \edb_top_inst/n2831 , 
        \edb_top_inst/n2832 , \edb_top_inst/n2833 , \edb_top_inst/n2834 , 
        \edb_top_inst/n2835 , \edb_top_inst/n2836 , \edb_top_inst/n2837 , 
        \edb_top_inst/n2838 , \edb_top_inst/n2839 , \edb_top_inst/n2840 , 
        \edb_top_inst/n2841 , \edb_top_inst/n2842 , \edb_top_inst/n2843 , 
        \edb_top_inst/n2844 , \edb_top_inst/n2845 , \edb_top_inst/n2846 , 
        \edb_top_inst/n2847 , \edb_top_inst/n2848 , \edb_top_inst/n2849 , 
        \edb_top_inst/n2850 , \edb_top_inst/n2851 , \edb_top_inst/n2852 , 
        \edb_top_inst/n2853 , \edb_top_inst/n2854 , \edb_top_inst/n2855 , 
        \edb_top_inst/n2856 , \edb_top_inst/n2857 , \edb_top_inst/n2858 , 
        \edb_top_inst/n2859 , \edb_top_inst/n2860 , \edb_top_inst/n2861 , 
        \edb_top_inst/n2862 , \edb_top_inst/n2863 , \edb_top_inst/n2864 , 
        \edb_top_inst/n2865 , \edb_top_inst/n2866 , \edb_top_inst/n2867 , 
        \edb_top_inst/n2868 , \edb_top_inst/n2869 , \edb_top_inst/n2870 , 
        \edb_top_inst/n2871 , \edb_top_inst/n2872 , \edb_top_inst/n2873 , 
        \edb_top_inst/n2874 , \edb_top_inst/n2875 , \edb_top_inst/n2876 , 
        \edb_top_inst/n2877 , \edb_top_inst/n2878 , \edb_top_inst/n2879 , 
        \edb_top_inst/n2880 , \edb_top_inst/n2881 , \edb_top_inst/n2882 , 
        \edb_top_inst/n2888 , \edb_top_inst/n2889 , \edb_top_inst/n2890 , 
        \edb_top_inst/n2891 , \edb_top_inst/n2892 , \edb_top_inst/n2893 , 
        \edb_top_inst/n2894 , \edb_top_inst/n2895 , \edb_top_inst/n2896 , 
        \edb_top_inst/n2897 , \edb_top_inst/n2898 , \edb_top_inst/n2899 , 
        \edb_top_inst/n2900 , \edb_top_inst/n2901 , \edb_top_inst/n2902 , 
        \edb_top_inst/n2903 , \edb_top_inst/n2904 , \edb_top_inst/n2905 , 
        \edb_top_inst/n2906 , \edb_top_inst/n2907 , \edb_top_inst/n2908 , 
        \edb_top_inst/n2909 , \edb_top_inst/n2910 , \edb_top_inst/n2911 , 
        \edb_top_inst/n2912 , \edb_top_inst/n2913 , \edb_top_inst/n2914 , 
        \edb_top_inst/n2915 , \edb_top_inst/n2916 , \edb_top_inst/n2917 , 
        \edb_top_inst/n2918 , \edb_top_inst/n2919 , \edb_top_inst/n2920 , 
        \edb_top_inst/n2921 , \edb_top_inst/n2922 , \edb_top_inst/n2923 , 
        \edb_top_inst/n2924 , \edb_top_inst/n2925 , \edb_top_inst/n2926 , 
        \edb_top_inst/n2927 , \edb_top_inst/n2928 , \edb_top_inst/n2929 , 
        \edb_top_inst/n2930 , \edb_top_inst/n2931 , \edb_top_inst/n2932 , 
        \edb_top_inst/n2933 , \edb_top_inst/n2934 , \edb_top_inst/n2935 , 
        \edb_top_inst/n2936 , \edb_top_inst/n2937 , \edb_top_inst/n2938 , 
        \edb_top_inst/n2939 , \edb_top_inst/n2940 , \edb_top_inst/n2941 , 
        \edb_top_inst/n2942 , \edb_top_inst/n2943 , \edb_top_inst/n2944 , 
        \edb_top_inst/n2945 , \edb_top_inst/n2946 , \edb_top_inst/n2947 , 
        \edb_top_inst/n2948 , \edb_top_inst/n2949 , \edb_top_inst/n2950 , 
        \edb_top_inst/n2951 , \edb_top_inst/n2952 , \edb_top_inst/n2953 , 
        \edb_top_inst/n2954 , \edb_top_inst/n2955 , \edb_top_inst/n2956 , 
        \edb_top_inst/n2957 , \edb_top_inst/n2958 , \edb_top_inst/n2959 , 
        \edb_top_inst/n2960 , \edb_top_inst/n2961 , \edb_top_inst/n2962 , 
        \edb_top_inst/n2963 , \edb_top_inst/n2964 , \edb_top_inst/n2965 , 
        \edb_top_inst/n2966 , \edb_top_inst/n2967 , \edb_top_inst/n2968 , 
        \edb_top_inst/n2969 , \edb_top_inst/n2970 , \edb_top_inst/n2971 , 
        \edb_top_inst/n2972 , \edb_top_inst/n2973 , \edb_top_inst/n2974 , 
        \edb_top_inst/n2975 , \edb_top_inst/n2976 , \edb_top_inst/n2977 , 
        \edb_top_inst/n2978 , \edb_top_inst/n2979 , \edb_top_inst/n2980 , 
        \edb_top_inst/n2981 , \edb_top_inst/n2982 , \edb_top_inst/n2983 , 
        \edb_top_inst/n2984 , \edb_top_inst/n2985 , \edb_top_inst/n2986 , 
        \edb_top_inst/n2987 , \edb_top_inst/n2988 , \edb_top_inst/n2989 , 
        \edb_top_inst/n2990 , \edb_top_inst/n2991 , \edb_top_inst/n2992 , 
        \edb_top_inst/n2993 , \edb_top_inst/n2994 , \edb_top_inst/n2995 , 
        \edb_top_inst/n2996 , \edb_top_inst/n2997 , \edb_top_inst/n2998 , 
        \edb_top_inst/n2999 , \edb_top_inst/n3000 , \edb_top_inst/n3001 , 
        \edb_top_inst/n3002 , \edb_top_inst/n3003 , \edb_top_inst/n3004 , 
        \edb_top_inst/n3005 , \edb_top_inst/n3006 , \edb_top_inst/n3007 , 
        \edb_top_inst/n3008 , \edb_top_inst/n3009 , \edb_top_inst/n3010 , 
        \edb_top_inst/n3011 , \edb_top_inst/n3012 , \edb_top_inst/n3013 , 
        \edb_top_inst/n3014 , \edb_top_inst/n3015 , \edb_top_inst/n3016 , 
        \edb_top_inst/n3017 , \edb_top_inst/n3018 , \edb_top_inst/n3019 , 
        \edb_top_inst/n3020 , \edb_top_inst/n3021 , \edb_top_inst/n3022 , 
        \edb_top_inst/n3023 , \edb_top_inst/n3024 , \edb_top_inst/n3025 , 
        \edb_top_inst/n3026 , \edb_top_inst/n3027 , \edb_top_inst/n3028 , 
        \edb_top_inst/n3029 , \edb_top_inst/n3030 , \edb_top_inst/n3031 , 
        \edb_top_inst/n3032 , \edb_top_inst/n3033 , \edb_top_inst/n3034 , 
        \edb_top_inst/n3035 , \edb_top_inst/n3036 , \edb_top_inst/n3037 , 
        \edb_top_inst/n3038 , \edb_top_inst/n3039 , \edb_top_inst/n3040 , 
        \edb_top_inst/n3041 , \edb_top_inst/n3042 , \edb_top_inst/n3043 , 
        \edb_top_inst/n3044 , \edb_top_inst/n3045 , \edb_top_inst/n3046 , 
        \edb_top_inst/n3047 , \edb_top_inst/n3048 , \edb_top_inst/n3049 , 
        \edb_top_inst/n3050 , \edb_top_inst/n3051 , \edb_top_inst/n3052 , 
        \edb_top_inst/n3053 , \edb_top_inst/n3054 , \edb_top_inst/n3055 , 
        \edb_top_inst/n3056 , \edb_top_inst/n3057 , \edb_top_inst/n3058 , 
        \edb_top_inst/n3059 , \edb_top_inst/n3060 , \edb_top_inst/n3061 , 
        \edb_top_inst/n3062 , \edb_top_inst/n3063 , \edb_top_inst/n3064 , 
        \edb_top_inst/n3065 , \edb_top_inst/n3066 , \edb_top_inst/n3067 , 
        \edb_top_inst/n3068 , \edb_top_inst/n3069 , \edb_top_inst/n3070 , 
        \edb_top_inst/n3071 , \edb_top_inst/n3072 , \edb_top_inst/n3073 , 
        \edb_top_inst/n3074 , \edb_top_inst/n3075 , \edb_top_inst/n3076 , 
        \edb_top_inst/n3077 , \edb_top_inst/n3078 , \edb_top_inst/n3079 , 
        \edb_top_inst/n3080 , \edb_top_inst/n3081 , \edb_top_inst/n3082 , 
        \edb_top_inst/n3083 , \edb_top_inst/n3084 , \edb_top_inst/n3085 , 
        \edb_top_inst/n3086 , \edb_top_inst/n3087 , \edb_top_inst/n3088 , 
        \edb_top_inst/n3089 , \edb_top_inst/n3090 , \edb_top_inst/n3091 , 
        \edb_top_inst/n3092 , \edb_top_inst/n3093 , \edb_top_inst/n3094 , 
        \edb_top_inst/n3095 , \edb_top_inst/n3096 , \edb_top_inst/n3097 , 
        \edb_top_inst/n3098 , \edb_top_inst/n3099 , \edb_top_inst/n3100 , 
        \edb_top_inst/n3101 , \edb_top_inst/n3102 , \edb_top_inst/n3103 , 
        \edb_top_inst/n3104 , \edb_top_inst/n3105 , \edb_top_inst/n3106 , 
        \edb_top_inst/n3107 , \edb_top_inst/n3108 , \edb_top_inst/n3109 , 
        \edb_top_inst/n3110 , \edb_top_inst/n3111 , \edb_top_inst/n3112 , 
        \edb_top_inst/n3113 , \edb_top_inst/n3114 , \edb_top_inst/n3115 , 
        \edb_top_inst/n3116 , \edb_top_inst/n3117 , \edb_top_inst/n3118 , 
        \edb_top_inst/n3119 , \edb_top_inst/n3120 , \edb_top_inst/n3121 , 
        \edb_top_inst/n3122 , \edb_top_inst/n3123 , \edb_top_inst/n3124 , 
        \edb_top_inst/n3125 , \edb_top_inst/n3126 , \edb_top_inst/n3127 , 
        \edb_top_inst/n3128 , \edb_top_inst/n3129 , \edb_top_inst/n3130 , 
        \edb_top_inst/n3131 , \edb_top_inst/n3132 , \edb_top_inst/n3133 , 
        \edb_top_inst/n3134 , \edb_top_inst/n3135 , \edb_top_inst/n3136 , 
        \edb_top_inst/n3137 , \edb_top_inst/n3138 , \edb_top_inst/n3139 , 
        \edb_top_inst/n3140 , \edb_top_inst/n3141 , \edb_top_inst/n3142 , 
        \edb_top_inst/n3143 , \edb_top_inst/n3144 , \edb_top_inst/n3145 , 
        \edb_top_inst/n3146 , \edb_top_inst/n3147 , \edb_top_inst/n3148 , 
        \edb_top_inst/n3149 , \edb_top_inst/n3150 , \edb_top_inst/n3151 , 
        \edb_top_inst/n3152 , \edb_top_inst/n3153 , \edb_top_inst/n3154 , 
        \edb_top_inst/n3155 , \edb_top_inst/n3156 , \edb_top_inst/n3157 , 
        \edb_top_inst/n3158 , \edb_top_inst/n3159 , \edb_top_inst/n3160 , 
        \edb_top_inst/n3161 , \edb_top_inst/n3162 , \edb_top_inst/n3163 , 
        \edb_top_inst/n3164 , \edb_top_inst/n3165 , \edb_top_inst/n3166 , 
        \edb_top_inst/n3167 , \edb_top_inst/n3168 , \edb_top_inst/n3169 , 
        \edb_top_inst/n3170 , \edb_top_inst/n3171 , \edb_top_inst/n3172 , 
        \edb_top_inst/n3173 , \edb_top_inst/n3174 , \edb_top_inst/n3175 , 
        \edb_top_inst/n3176 , \edb_top_inst/n3177 , \edb_top_inst/n3178 , 
        \edb_top_inst/n3179 , \edb_top_inst/n3180 , \edb_top_inst/n3181 , 
        \edb_top_inst/n3182 , \edb_top_inst/n3183 , \edb_top_inst/n3184 , 
        \edb_top_inst/n3185 , \edb_top_inst/n3186 , \edb_top_inst/n3187 , 
        \edb_top_inst/n3188 , \edb_top_inst/n3189 , \edb_top_inst/n3190 , 
        \edb_top_inst/n3191 , \edb_top_inst/n3192 , \edb_top_inst/n3193 , 
        \edb_top_inst/n3194 , \edb_top_inst/n3195 , \edb_top_inst/n3196 , 
        \edb_top_inst/n3197 , \edb_top_inst/n3198 , \edb_top_inst/n3199 , 
        \edb_top_inst/n3200 , \edb_top_inst/n3201 , \edb_top_inst/n3202 , 
        \edb_top_inst/n3203 , \edb_top_inst/n3204 , \edb_top_inst/n3205 , 
        \edb_top_inst/n3206 , \edb_top_inst/n3207 , \edb_top_inst/n3208 , 
        \edb_top_inst/n3209 , \edb_top_inst/n3210 , \edb_top_inst/n3211 , 
        \edb_top_inst/n3212 , \edb_top_inst/n3213 , \edb_top_inst/n3214 , 
        \edb_top_inst/n3215 , \edb_top_inst/n3216 , \edb_top_inst/n3217 , 
        \edb_top_inst/n3218 , \edb_top_inst/n3219 , \edb_top_inst/n3220 , 
        \edb_top_inst/n3221 , \edb_top_inst/n3222 , \edb_top_inst/n3223 , 
        \edb_top_inst/n3224 , \edb_top_inst/n3225 , \edb_top_inst/n3226 , 
        \edb_top_inst/n3227 , \edb_top_inst/n3228 , \edb_top_inst/n3229 , 
        \edb_top_inst/n3230 , \edb_top_inst/n3231 , \edb_top_inst/n3232 , 
        \edb_top_inst/n3233 , \edb_top_inst/n3234 , \edb_top_inst/n3235 , 
        \edb_top_inst/n3236 , \edb_top_inst/n3237 , \edb_top_inst/n3238 , 
        \edb_top_inst/n3239 , \edb_top_inst/n3240 , \edb_top_inst/n3241 , 
        \edb_top_inst/n3242 , \edb_top_inst/n3243 , \edb_top_inst/n3244 , 
        \edb_top_inst/n3245 , \edb_top_inst/n3246 , \edb_top_inst/n3247 , 
        \edb_top_inst/n3248 , \edb_top_inst/n3249 , \edb_top_inst/n3250 , 
        \edb_top_inst/n3251 , \edb_top_inst/n3252 , \edb_top_inst/n3253 , 
        \edb_top_inst/n3254 , \edb_top_inst/n3255 , \edb_top_inst/n3256 , 
        \edb_top_inst/n3257 , \edb_top_inst/n3258 , \edb_top_inst/n3259 , 
        \edb_top_inst/n3260 , \edb_top_inst/n3261 , \edb_top_inst/n3262 , 
        \edb_top_inst/n3263 , \edb_top_inst/n3264 , \edb_top_inst/n3265 , 
        \edb_top_inst/n3266 , \edb_top_inst/n3267 , \edb_top_inst/n3268 , 
        \edb_top_inst/n3269 , \edb_top_inst/n3270 , \edb_top_inst/n3271 , 
        \edb_top_inst/n3272 , \edb_top_inst/n3273 , \edb_top_inst/n3274 , 
        \edb_top_inst/n3275 , \edb_top_inst/n3276 , \edb_top_inst/n3277 , 
        \edb_top_inst/n3278 , \edb_top_inst/n3279 , \edb_top_inst/n3280 , 
        \edb_top_inst/n3281 , \edb_top_inst/n3282 , \edb_top_inst/n3283 , 
        \edb_top_inst/n3284 , \edb_top_inst/n3285 , \edb_top_inst/n3286 , 
        \edb_top_inst/n3287 , \edb_top_inst/n3288 , \edb_top_inst/n3289 , 
        \edb_top_inst/n3290 , \edb_top_inst/n3291 , \edb_top_inst/n3292 , 
        \edb_top_inst/n3293 , \edb_top_inst/n3294 , \edb_top_inst/n3295 , 
        \edb_top_inst/n3296 , \edb_top_inst/n3297 , \edb_top_inst/n3298 , 
        \edb_top_inst/n3299 , \edb_top_inst/n3300 , \edb_top_inst/n3301 , 
        \edb_top_inst/n3302 , \edb_top_inst/n3303 , \edb_top_inst/n3304 , 
        \edb_top_inst/n3305 , \edb_top_inst/n3306 , \edb_top_inst/n3307 , 
        \edb_top_inst/n3308 , \edb_top_inst/n3309 , \edb_top_inst/n3310 , 
        \edb_top_inst/n3311 , \edb_top_inst/n3312 , \edb_top_inst/n3313 , 
        \edb_top_inst/n3314 , \edb_top_inst/n3315 , \edb_top_inst/n3316 , 
        \edb_top_inst/n3317 , \edb_top_inst/n3318 , \edb_top_inst/n3319 , 
        \edb_top_inst/n3320 , \edb_top_inst/n3321 , \edb_top_inst/n3322 , 
        \edb_top_inst/n3323 , \edb_top_inst/n3324 , \edb_top_inst/n3325 , 
        \edb_top_inst/n3326 , \edb_top_inst/n3327 , \edb_top_inst/n3328 , 
        \edb_top_inst/n3329 , \edb_top_inst/n3330 , \edb_top_inst/n3331 , 
        \edb_top_inst/n3332 , \edb_top_inst/n3333 , \edb_top_inst/n3334 , 
        \edb_top_inst/n3335 , \edb_top_inst/n3336 , \edb_top_inst/n3337 , 
        \edb_top_inst/n3338 , \edb_top_inst/n3339 , \edb_top_inst/n3340 , 
        \edb_top_inst/n2739 , n3357, n3358, n3359, n3360, n3361, 
        n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, 
        n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, 
        n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, 
        n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, 
        n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, 
        n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, 
        n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, 
        n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, 
        n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, 
        n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, 
        n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, 
        n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, 
        n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, 
        n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, 
        n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, 
        n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, 
        n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, 
        n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, 
        n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, 
        n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, 
        n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, 
        n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, 
        n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, 
        n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, 
        n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, 
        n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, 
        n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, 
        n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, 
        n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, 
        n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, 
        n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, 
        n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, 
        n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, 
        n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, 
        n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, 
        n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, 
        n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, 
        n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, 
        n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, 
        n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, 
        n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, 
        n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, 
        n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, 
        n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, 
        n3714, n3715, n3716, n3717, n3718, n3726, n3727, n3728, 
        n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, 
        n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, 
        n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, 
        n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, 
        n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, 
        n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, 
        n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, 
        n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, 
        n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, 
        n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, 
        n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, 
        n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, 
        n3825, n3826, n3827, n3828, n3829, wCdcFifoFull, rSRST, 
        \MCsiRxController/n279 , \MCsiRxController/MCsi2Decoder/n630 , \MCsiRxController/MCsi2Decoder/n632 , 
        \MCsiRxController/MCsi2Decoder/n7 , \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[0] , \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRVd , 
        \~MCsiRxController/MCsi2Decoder/reduce_nor_75/n1 , \MCsiRxController/MCsi2Decoder/n603 , 
        \MCsiRxController/MCsi2Decoder/qLineCntRst , \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE , 
        \MCsiRxController/MCsi2Decoder/n96 , \MCsiRxController/MCsi2Decoder/n606 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/equal_38/n19 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n233 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n238 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n243 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n248 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n253 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n258 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n263 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n268 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n273 , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[1] , \MCsiRxController/MCsi2Decoder/wFtiRd[2] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[3] , \MCsiRxController/MCsi2Decoder/wFtiRd[4] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[5] , \MCsiRxController/MCsi2Decoder/wFtiRd[6] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[7] , \MCsiRxController/MCsi2Decoder/wFtiRd[8] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[9] , \MCsiRxController/MCsi2Decoder/wFtiRd[10] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[11] , \MCsiRxController/MCsi2Decoder/wFtiRd[12] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[13] , \MCsiRxController/MCsi2Decoder/wFtiRd[14] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[15] , \MCsiRxController/MCsi2Decoder/equal_62/n5 , 
        \MCsiRxController/MCsi2Decoder/equal_59/n5 , \MCsiRxController/genblk1[0].mVideoFIFO/qRE , 
        \MCsiRxController/genblk1[0].mVideoFIFO/qFullAllmost , \MCsiRxController/genblk1[0].mVideoFIFO/qRVD , 
        \MCsiRxController/genblk1[0].mVideoFIFO/equal_75/n17 , \MCsiRxController/genblk1[0].mVideoFIFO/n436 , 
        \MCsiRxController/genblk1[0].mVideoFIFO/n441 , \MCsiRxController/genblk1[0].mVideoFIFO/n446 , 
        \MCsiRxController/genblk1[0].mVideoFIFO/n451 , \MCsiRxController/genblk1[0].mVideoFIFO/n456 , 
        \MCsiRxController/genblk1[0].mVideoFIFO/n461 , \MCsiRxController/genblk1[0].mVideoFIFO/n466 , 
        \MCsiRxController/genblk1[0].mVideoFIFO/n471 , \MCsiRxController/n278 , 
        \MCsiRxController/n277 , \MCsiRxController/n276 , \MCsiRxController/n275 , 
        \MCsiRxController/n274 , \MCsiRxController/n273 , \MCsiRxController/n272 , 
        \MCsiRxController/n271 , \MCsiRxController/n270 , \MCsiRxController/n269 , 
        \MCsiRxController/n268 , \MCsiRxController/n267 , \MCsiRxController/n266 , 
        \MCsiRxController/n265 , \MCsiRxController/n264 , \MVideoPostProcess/qVtgRstCntCke , 
        \MVideoPostProcess/rVtgRstSel , \MVideoPostProcess/equal_18/n21 , 
        \~n1834 , ceg_net939, \MVideoPostProcess/inst_adv7511_config/n816 , 
        \MVideoPostProcess/inst_adv7511_config/n833 , \~ceg_net512 , \MVideoPostProcess/inst_adv7511_config/n268 , 
        ceg_net995, \MVideoPostProcess/inst_adv7511_config/n1107 , \MVideoPostProcess/inst_adv7511_config/n1224 , 
        \MVideoPostProcess/inst_adv7511_config/n277 , ceg_net479, \MVideoPostProcess/inst_adv7511_config/n242 , 
        ceg_net1327, \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15] , 
        \MVideoPostProcess/inst_adv7511_config/n1243 , \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n846 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n852 , 
        ceg_net1087, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n847 , 
        ceg_net1335, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n848 , 
        ceg_net566, \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] , 
        ceg_net1400, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n870 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n879 , 
        ceg_net1463, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n829 , 
        ceg_net1361, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n899 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n898 , 
        ceg_net616, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n845 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n844 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n843 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n842 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n841 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n840 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n839 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n851 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n850 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n869 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n868 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n867 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n866 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n865 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n864 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n863 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n878 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n877 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n876 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n875 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n874 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n873 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n872 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n828 , 
        ceg_net1471, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n827 , 
        ceg_net1480, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n826 , 
        ceg_net1488, n10139, n10138, n10137, n10136, \MVideoPostProcess/mVideoTimingGen/qVrange , 
        \MVideoPostProcess/rVtgRST[2] , \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2 , 
        \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1 , \MVideoPostProcess/inst_adv7511_config/n251 , 
        \MVideoPostProcess/inst_adv7511_config/n250 , \MVideoPostProcess/inst_adv7511_config/n249 , 
        \MVideoPostProcess/inst_adv7511_config/n248 , \MVideoPostProcess/inst_adv7511_config/n247 , 
        \MVideoPostProcess/inst_adv7511_config/n246 , \MVideoPostProcess/inst_adv7511_config/n245 , 
        \MVideoPostProcess/inst_adv7511_config/n244 , \MVideoPostProcess/inst_adv7511_config/n700 , 
        \MVideoPostProcess/inst_adv7511_config/n705 , \MVideoPostProcess/inst_adv7511_config/n710 , 
        \MVideoPostProcess/inst_adv7511_config/n715 , \MVideoPostProcess/inst_adv7511_config/n720 , 
        \MVideoPostProcess/inst_adv7511_config/n725 , \MVideoPostProcess/inst_adv7511_config/n730 , 
        \MVideoPostProcess/inst_adv7511_config/n735 , \MVideoPostProcess/inst_adv7511_config/n740 , 
        \MVideoPostProcess/inst_adv7511_config/n745 , \MVideoPostProcess/inst_adv7511_config/n750 , 
        \MVideoPostProcess/inst_adv7511_config/n755 , \MVideoPostProcess/inst_adv7511_config/n760 , 
        \MVideoPostProcess/inst_adv7511_config/n765 , \MVideoPostProcess/inst_adv7511_config/n770 , 
        \MVideoPostProcess/inst_adv7511_config/n780 , \MVideoPostProcess/inst_adv7511_config/n785 , 
        \MVideoPostProcess/inst_adv7511_config/n790 , \MVideoPostProcess/inst_adv7511_config/n795 , 
        \MVideoPostProcess/inst_adv7511_config/n800 , \MVideoPostProcess/inst_adv7511_config/n805 , 
        \MVideoPostProcess/inst_adv7511_config/n810 , \MVideoPostProcess/inst_adv7511_config/n276 , 
        \MVideoPostProcess/inst_adv7511_config/n275 , \MVideoPostProcess/inst_adv7511_config/n274 , 
        \MVideoPostProcess/inst_adv7511_config/n273 , \MVideoPostProcess/inst_adv7511_config/n272 , 
        \MVideoPostProcess/inst_adv7511_config/n271 , \MVideoPostProcess/inst_adv7511_config/n270 , 
        \MVideoPostProcess/mVideoTimingGen/n131 , \MVideoPostProcess/mVideoTimingGen/equal_12/n23 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] , 
        \MVideoPostProcess/mVideoTimingGen/qVde , \MVideoPostProcess/mVideoTimingGen/n267 , 
        \MVideoPostProcess/mVideoTimingGen/rHSync[3] , \MVideoPostProcess/mVideoTimingGen/n130 , 
        \MVideoPostProcess/mVideoTimingGen/n129 , \MVideoPostProcess/mVideoTimingGen/n126 , 
        \MVideoPostProcess/mVideoTimingGen/n125 , \MVideoPostProcess/mVideoTimingGen/n121 , 
        \MVideoPostProcess/mVideoTimingGen/qHrange , \MVideoPostProcess/mVideoTimingGen/rVSync[3] , 
        \MVideoPostProcess/wVgaGenFDe , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qFullAllmost , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n478 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n483 , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n488 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n493 , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n498 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n503 , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n508 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n513 , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n518 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n523 , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n528 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n533 , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12] , 
        \genblk1.genblk1[0].mPulseGenerator/equal_6/n5 , \genblk1.genblk1[0].mPulseGenerator/equal_12/n25 , 
        \genblk1.genblk1[3].mPulseGenerator/equal_6/n5 , \genblk1.genblk1[3].mPulseGenerator/n50 , 
        \genblk1.genblk1[4].mPulseGenerator/equal_6/n5 , \genblk1.genblk1[4].mPulseGenerator/n50 , 
        \edb_top_inst/la0/n1340 , \edb_top_inst/ceg_net5 , \edb_top_inst/edb_user_dr[60] , 
        \edb_top_inst/la0/n1312 , \edb_top_inst/la0/n1341 , \edb_top_inst/la0/n1342 , 
        \edb_top_inst/edb_user_dr[62] , \edb_top_inst/edb_user_dr[0] , \edb_top_inst/la0/n1396 , 
        \edb_top_inst/edb_user_dr[42] , \edb_top_inst/la0/n1913 , \edb_top_inst/edb_user_dr[59] , 
        \edb_top_inst/la0/n1965 , \edb_top_inst/la0/data_to_addr_counter[0] , 
        \edb_top_inst/la0/addr_ct_en , \edb_top_inst/edb_user_dr[77] , \edb_top_inst/la0/op_reg_en , 
        \edb_top_inst/la0/n2189 , \edb_top_inst/ceg_net26 , \edb_top_inst/la0/data_to_word_counter[0] , 
        \edb_top_inst/la0/word_ct_en , \edb_top_inst/la0/n2466 , \edb_top_inst/ceg_net14 , 
        \edb_top_inst/la0/module_next_state[0] , la0_probe1, \edb_top_inst/la0/n5294 , 
        \edb_top_inst/la0/n5492 , \edb_top_inst/la0/n6947 , \edb_top_inst/la0/n7907 , 
        \edb_top_inst/la0/n8105 , \edb_top_inst/la0/n8741 , \edb_top_inst/la0/n9645 , 
        \edb_top_inst/la0/n9843 , \edb_top_inst/la0/n10527 , \edb_top_inst/la0/n10542 , 
        \edb_top_inst/la0/n10740 , \edb_top_inst/la0/n11368 , \edb_top_inst/la0/n12201 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/edb_user_dr[64] , \edb_top_inst/la0/regsel_ld_en , 
        \edb_top_inst/edb_user_dr[43] , \edb_top_inst/edb_user_dr[61] , 
        \edb_top_inst/edb_user_dr[63] , \edb_top_inst/edb_user_dr[1] , \edb_top_inst/edb_user_dr[2] , 
        \edb_top_inst/edb_user_dr[3] , \edb_top_inst/edb_user_dr[4] , \edb_top_inst/edb_user_dr[5] , 
        \edb_top_inst/edb_user_dr[6] , \edb_top_inst/edb_user_dr[7] , \edb_top_inst/edb_user_dr[8] , 
        \edb_top_inst/edb_user_dr[9] , \edb_top_inst/edb_user_dr[10] , \edb_top_inst/edb_user_dr[11] , 
        \edb_top_inst/edb_user_dr[12] , \edb_top_inst/edb_user_dr[13] , 
        \edb_top_inst/edb_user_dr[14] , \edb_top_inst/edb_user_dr[15] , 
        \edb_top_inst/edb_user_dr[16] , \edb_top_inst/edb_user_dr[17] , 
        \edb_top_inst/edb_user_dr[18] , \edb_top_inst/edb_user_dr[19] , 
        \edb_top_inst/edb_user_dr[20] , \edb_top_inst/edb_user_dr[21] , 
        \edb_top_inst/edb_user_dr[22] , \edb_top_inst/edb_user_dr[23] , 
        \edb_top_inst/edb_user_dr[24] , \edb_top_inst/edb_user_dr[25] , 
        \edb_top_inst/edb_user_dr[26] , \edb_top_inst/edb_user_dr[27] , 
        \edb_top_inst/edb_user_dr[28] , \edb_top_inst/edb_user_dr[29] , 
        \edb_top_inst/edb_user_dr[30] , \edb_top_inst/edb_user_dr[31] , 
        \edb_top_inst/edb_user_dr[32] , \edb_top_inst/edb_user_dr[33] , 
        \edb_top_inst/edb_user_dr[34] , \edb_top_inst/edb_user_dr[35] , 
        \edb_top_inst/edb_user_dr[36] , \edb_top_inst/edb_user_dr[37] , 
        \edb_top_inst/edb_user_dr[38] , \edb_top_inst/edb_user_dr[39] , 
        \edb_top_inst/edb_user_dr[40] , \edb_top_inst/edb_user_dr[41] , 
        \edb_top_inst/edb_user_dr[44] , \edb_top_inst/edb_user_dr[45] , 
        \edb_top_inst/edb_user_dr[46] , \edb_top_inst/edb_user_dr[47] , 
        \edb_top_inst/edb_user_dr[48] , \edb_top_inst/edb_user_dr[49] , 
        \edb_top_inst/edb_user_dr[50] , \edb_top_inst/edb_user_dr[51] , 
        \edb_top_inst/edb_user_dr[52] , \edb_top_inst/edb_user_dr[53] , 
        \edb_top_inst/edb_user_dr[54] , \edb_top_inst/edb_user_dr[55] , 
        \edb_top_inst/edb_user_dr[56] , \edb_top_inst/edb_user_dr[57] , 
        \edb_top_inst/edb_user_dr[58] , \edb_top_inst/la0/data_to_addr_counter[1] , 
        \edb_top_inst/la0/data_to_addr_counter[2] , \edb_top_inst/la0/data_to_addr_counter[3] , 
        \edb_top_inst/la0/data_to_addr_counter[4] , \edb_top_inst/la0/data_to_addr_counter[5] , 
        \edb_top_inst/la0/data_to_addr_counter[6] , \edb_top_inst/la0/data_to_addr_counter[7] , 
        \edb_top_inst/la0/data_to_addr_counter[8] , \edb_top_inst/la0/data_to_addr_counter[9] , 
        \edb_top_inst/la0/data_to_addr_counter[10] , \edb_top_inst/la0/data_to_addr_counter[11] , 
        \edb_top_inst/la0/data_to_addr_counter[12] , \edb_top_inst/la0/data_to_addr_counter[13] , 
        \edb_top_inst/la0/data_to_addr_counter[14] , \edb_top_inst/la0/data_to_addr_counter[15] , 
        \edb_top_inst/la0/data_to_addr_counter[16] , \edb_top_inst/la0/data_to_addr_counter[17] , 
        \edb_top_inst/la0/data_to_addr_counter[18] , \edb_top_inst/la0/data_to_addr_counter[19] , 
        \edb_top_inst/la0/data_to_addr_counter[20] , \edb_top_inst/la0/data_to_addr_counter[21] , 
        \edb_top_inst/la0/data_to_addr_counter[22] , \edb_top_inst/la0/data_to_addr_counter[23] , 
        \edb_top_inst/la0/data_to_addr_counter[24] , \edb_top_inst/la0/data_to_addr_counter[25] , 
        \edb_top_inst/la0/data_to_addr_counter[26] , \edb_top_inst/edb_user_dr[78] , 
        \edb_top_inst/edb_user_dr[79] , \edb_top_inst/edb_user_dr[80] , 
        \edb_top_inst/la0/n2188 , \edb_top_inst/la0/n2187 , \edb_top_inst/la0/n2186 , 
        \edb_top_inst/la0/n2185 , \edb_top_inst/la0/n2184 , \edb_top_inst/la0/data_to_word_counter[1] , 
        \edb_top_inst/la0/data_to_word_counter[2] , \edb_top_inst/la0/data_to_word_counter[3] , 
        \edb_top_inst/la0/data_to_word_counter[4] , \edb_top_inst/la0/data_to_word_counter[5] , 
        \edb_top_inst/la0/data_to_word_counter[6] , \edb_top_inst/la0/data_to_word_counter[7] , 
        \edb_top_inst/la0/data_to_word_counter[8] , \edb_top_inst/la0/data_to_word_counter[9] , 
        \edb_top_inst/la0/data_to_word_counter[10] , \edb_top_inst/la0/data_to_word_counter[11] , 
        \edb_top_inst/la0/data_to_word_counter[12] , \edb_top_inst/la0/data_to_word_counter[13] , 
        \edb_top_inst/la0/data_to_word_counter[14] , \edb_top_inst/la0/data_to_word_counter[15] , 
        \edb_top_inst/la0/n2465 , \edb_top_inst/la0/n2464 , \edb_top_inst/la0/n2463 , 
        \edb_top_inst/la0/n2462 , \edb_top_inst/la0/n2461 , \edb_top_inst/la0/n2460 , 
        \edb_top_inst/la0/n2459 , \edb_top_inst/la0/n2458 , \edb_top_inst/la0/n2457 , 
        \edb_top_inst/la0/n2456 , \edb_top_inst/la0/n2455 , \edb_top_inst/la0/n2454 , 
        \edb_top_inst/la0/n2453 , \edb_top_inst/la0/n2452 , \edb_top_inst/la0/n2451 , 
        \edb_top_inst/la0/n2450 , \edb_top_inst/la0/n2449 , \edb_top_inst/la0/n2448 , 
        \edb_top_inst/la0/n2447 , \edb_top_inst/la0/n2446 , \edb_top_inst/la0/n2445 , 
        \edb_top_inst/la0/n2444 , \edb_top_inst/la0/n2443 , \edb_top_inst/la0/n2442 , 
        \edb_top_inst/la0/n2441 , \edb_top_inst/la0/n2440 , \edb_top_inst/la0/n2439 , 
        \edb_top_inst/la0/n2438 , \edb_top_inst/la0/n2437 , \edb_top_inst/la0/n2436 , 
        \edb_top_inst/la0/n2435 , \edb_top_inst/la0/n2434 , \edb_top_inst/la0/n2433 , 
        \edb_top_inst/la0/n2432 , \edb_top_inst/la0/n2431 , \edb_top_inst/la0/n2430 , 
        \edb_top_inst/la0/n2429 , \edb_top_inst/la0/n2428 , \edb_top_inst/la0/n2427 , 
        \edb_top_inst/la0/n2426 , \edb_top_inst/la0/n2425 , \edb_top_inst/la0/n2424 , 
        \edb_top_inst/la0/n2423 , \edb_top_inst/la0/n2422 , \edb_top_inst/la0/n2421 , 
        \edb_top_inst/la0/n2420 , \edb_top_inst/la0/n2419 , \edb_top_inst/la0/n2418 , 
        \edb_top_inst/la0/n2417 , \edb_top_inst/la0/n2416 , \edb_top_inst/la0/n2415 , 
        \edb_top_inst/la0/n2414 , \edb_top_inst/la0/n2413 , \edb_top_inst/la0/n2412 , 
        \edb_top_inst/la0/n2411 , \edb_top_inst/la0/n2410 , \edb_top_inst/la0/n2409 , 
        \edb_top_inst/la0/n2408 , \edb_top_inst/la0/n2407 , \edb_top_inst/la0/n2406 , 
        \edb_top_inst/la0/n2405 , \edb_top_inst/la0/n2404 , \edb_top_inst/la0/n2403 , 
        \edb_top_inst/la0/module_next_state[1] , \edb_top_inst/la0/module_next_state[2] , 
        \edb_top_inst/la0/module_next_state[3] , \edb_top_inst/la0/axi_crc_i/n150 , 
        \edb_top_inst/ceg_net221 , \edb_top_inst/la0/axi_crc_i/n149 , \edb_top_inst/la0/axi_crc_i/n148 , 
        \edb_top_inst/la0/axi_crc_i/n147 , \edb_top_inst/la0/axi_crc_i/n146 , 
        \edb_top_inst/la0/axi_crc_i/n145 , \edb_top_inst/la0/axi_crc_i/n144 , 
        \edb_top_inst/la0/axi_crc_i/n143 , \edb_top_inst/la0/axi_crc_i/n142 , 
        \edb_top_inst/la0/axi_crc_i/n141 , \edb_top_inst/la0/axi_crc_i/n140 , 
        \edb_top_inst/la0/axi_crc_i/n139 , \edb_top_inst/la0/axi_crc_i/n138 , 
        \edb_top_inst/la0/axi_crc_i/n137 , \edb_top_inst/la0/axi_crc_i/n136 , 
        \edb_top_inst/la0/axi_crc_i/n135 , \edb_top_inst/la0/axi_crc_i/n134 , 
        \edb_top_inst/la0/axi_crc_i/n133 , \edb_top_inst/la0/axi_crc_i/n132 , 
        \edb_top_inst/la0/axi_crc_i/n131 , \edb_top_inst/la0/axi_crc_i/n130 , 
        \edb_top_inst/la0/axi_crc_i/n129 , \edb_top_inst/la0/axi_crc_i/n128 , 
        \edb_top_inst/la0/axi_crc_i/n127 , \edb_top_inst/la0/axi_crc_i/n126 , 
        \edb_top_inst/la0/axi_crc_i/n125 , \edb_top_inst/la0/axi_crc_i/n124 , 
        \edb_top_inst/la0/axi_crc_i/n123 , \edb_top_inst/la0/axi_crc_i/n122 , 
        \edb_top_inst/la0/axi_crc_i/n121 , \edb_top_inst/la0/axi_crc_i/n120 , 
        \edb_top_inst/la0/axi_crc_i/n119 , \edb_top_inst/la0/n2766 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/n3599 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/n4432 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/n5279 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n16 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n10 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n17 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/equal_9/n3 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n26 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n15 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n9 , \edb_top_inst/la0/n6114 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/n7892 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n72 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n38 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n73 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/equal_9/n31 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n82 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n71 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n70 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n69 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n68 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n67 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n66 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n65 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n64 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n63 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n62 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n61 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n60 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n59 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n58 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n57 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n37 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n36 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n35 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n34 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n33 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n32 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n31 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n30 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n29 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n28 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n27 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n26 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n25 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n24 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/n9630 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n40 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/equal_9/n15 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n50 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n39 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n38 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n37 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n36 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n35 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n34 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n33 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n21 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n20 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n19 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n18 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n17 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n16 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n15 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n22 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n41 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/equal_9/n15 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n50 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n39 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n38 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n37 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n36 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n35 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n34 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n33 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n21 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n19 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n18 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n17 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n16 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n15 , \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/trigger_tu/n89 , 
        \edb_top_inst/la0/la_biu_inst/next_state[0] , \edb_top_inst/la0/la_biu_inst/run_trig_p1 , 
        \edb_top_inst/la0/la_biu_inst/n382 , \edb_top_inst/la0/la_biu_inst/n1315 , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[0] , \edb_top_inst/la0/la_biu_inst/next_fsm_state[0] , 
        \edb_top_inst/ceg_net351 , \edb_top_inst/la0/la_biu_inst/n1300 , 
        \edb_top_inst/la0/n17781 , \edb_top_inst/la0/la_biu_inst/next_state[2] , 
        \edb_top_inst/la0/la_biu_inst/next_state[1] , \edb_top_inst/ceg_net348 , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[1] , \edb_top_inst/la0/la_biu_inst/fifo_dout[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[3] , \edb_top_inst/la0/la_biu_inst/fifo_dout[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[5] , \edb_top_inst/la0/la_biu_inst/fifo_dout[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[7] , \edb_top_inst/la0/la_biu_inst/fifo_dout[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[9] , \edb_top_inst/la0/la_biu_inst/fifo_dout[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[11] , \edb_top_inst/la0/la_biu_inst/fifo_dout[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[13] , \edb_top_inst/la0/la_biu_inst/fifo_dout[14] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[15] , \edb_top_inst/la0/la_biu_inst/fifo_dout[16] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[17] , \edb_top_inst/la0/la_biu_inst/fifo_dout[18] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[19] , \edb_top_inst/la0/la_biu_inst/fifo_dout[20] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[21] , \edb_top_inst/la0/la_biu_inst/fifo_dout[22] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[23] , \edb_top_inst/la0/la_biu_inst/fifo_dout[24] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[25] , \edb_top_inst/la0/la_biu_inst/fifo_dout[26] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[27] , \edb_top_inst/la0/la_biu_inst/fifo_dout[28] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[29] , \edb_top_inst/la0/la_biu_inst/fifo_dout[30] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[31] , \edb_top_inst/la0/la_biu_inst/fifo_dout[32] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[33] , \edb_top_inst/la0/la_biu_inst/fifo_dout[34] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[35] , \edb_top_inst/la0/la_biu_inst/fifo_dout[36] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[37] , \edb_top_inst/la0/la_biu_inst/fifo_dout[38] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[39] , \edb_top_inst/la0/la_biu_inst/fifo_dout[40] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[41] , \edb_top_inst/la0/la_biu_inst/fifo_dout[42] , 
        \edb_top_inst/la0/la_biu_inst/next_fsm_state[1] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data , 
        \edb_top_inst/la0/la_biu_inst/fifo_rstn , \edb_top_inst/la0/la_biu_inst/n2053 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 , \edb_top_inst/la0/la_biu_inst/fifo_push , 
        \edb_top_inst/ceg_net355 , \edb_top_inst/n73 , \edb_top_inst/n1044 , 
        \edb_top_inst/n1042 , \edb_top_inst/n1040 , \edb_top_inst/n1038 , 
        \edb_top_inst/n1036 , \edb_top_inst/n1034 , \edb_top_inst/n1032 , 
        \edb_top_inst/n1030 , \edb_top_inst/n1028 , \edb_top_inst/n1027 , 
        \edb_top_inst/n693 , \edb_top_inst/n1025 , \edb_top_inst/n1023 , 
        \edb_top_inst/n1021 , \edb_top_inst/n1019 , \edb_top_inst/n1017 , 
        \edb_top_inst/n1015 , \edb_top_inst/n1013 , \edb_top_inst/n1011 , 
        \edb_top_inst/n1008 , \edb_top_inst/n1005 , \edb_top_inst/n695 , 
        \edb_top_inst/n856 , \edb_top_inst/n854 , \edb_top_inst/n852 , 
        \edb_top_inst/n850 , \edb_top_inst/n848 , \edb_top_inst/n846 , 
        \edb_top_inst/n844 , \edb_top_inst/n842 , \edb_top_inst/n840 , 
        \edb_top_inst/n838 , \edb_top_inst/n710 , \edb_top_inst/n731 , 
        \edb_top_inst/n729 , \edb_top_inst/n727 , \edb_top_inst/n725 , 
        \edb_top_inst/n723 , \edb_top_inst/n721 , \edb_top_inst/n719 , 
        \edb_top_inst/n717 , \edb_top_inst/n715 , \edb_top_inst/n713 , 
        \edb_top_inst/n712 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[11] , 
        \edb_top_inst/n711 , \edb_top_inst/n752 , \edb_top_inst/n750 , 
        \edb_top_inst/n748 , \edb_top_inst/n746 , \edb_top_inst/n744 , 
        \edb_top_inst/n742 , \edb_top_inst/n740 , \edb_top_inst/n738 , 
        \edb_top_inst/n736 , \edb_top_inst/n734 , \edb_top_inst/n733 , 
        \edb_top_inst/edb_user_dr[65] , \edb_top_inst/edb_user_dr[66] , 
        \edb_top_inst/edb_user_dr[67] , \edb_top_inst/edb_user_dr[68] , 
        \edb_top_inst/edb_user_dr[69] , \edb_top_inst/edb_user_dr[70] , 
        \edb_top_inst/edb_user_dr[71] , \edb_top_inst/edb_user_dr[72] , 
        \edb_top_inst/edb_user_dr[73] , \edb_top_inst/edb_user_dr[74] , 
        \edb_top_inst/edb_user_dr[75] , \edb_top_inst/edb_user_dr[76] , 
        \edb_top_inst/debug_hub_inst/n266 , \edb_top_inst/debug_hub_inst/n95 , 
        \edb_top_inst/edb_user_dr[81] , \edb_top_inst/n714 , \edb_top_inst/n716 , 
        \edb_top_inst/n718 , \edb_top_inst/n720 , \edb_top_inst/n722 , 
        \edb_top_inst/n724 , \edb_top_inst/n726 , \edb_top_inst/n728 , 
        \edb_top_inst/n730 , \edb_top_inst/n732 , \edb_top_inst/n735 , 
        \edb_top_inst/n737 , \edb_top_inst/n739 , \edb_top_inst/n741 , 
        \edb_top_inst/n743 , \edb_top_inst/n745 , \edb_top_inst/n747 , 
        \edb_top_inst/n749 , \edb_top_inst/n751 , \edb_top_inst/n753 , 
        \edb_top_inst/n841 , \edb_top_inst/n843 , \edb_top_inst/n845 , 
        \edb_top_inst/n847 , \edb_top_inst/n849 , \edb_top_inst/n851 , 
        \edb_top_inst/n853 , \edb_top_inst/n855 , \edb_top_inst/n857 , 
        \edb_top_inst/n1009 , \edb_top_inst/n1012 , \edb_top_inst/n1014 , 
        \edb_top_inst/n1016 , \edb_top_inst/n1018 , \edb_top_inst/n1020 , 
        \edb_top_inst/n1022 , \edb_top_inst/n1024 , \edb_top_inst/n1026 , 
        \edb_top_inst/n1029 , \edb_top_inst/n1031 , \edb_top_inst/n1033 , 
        \edb_top_inst/n1035 , \edb_top_inst/n1037 , \edb_top_inst/n1039 , 
        \edb_top_inst/n1041 , \edb_top_inst/n1043 , \edb_top_inst/n1045 , 
        \edb_top_inst/n1048 , \edb_top_inst/n1050 , \edb_top_inst/n1052 , 
        \edb_top_inst/n1065 , \edb_top_inst/n1067 , \edb_top_inst/n1069 , 
        \edb_top_inst/n1071 , \edb_top_inst/n1073 , \edb_top_inst/n1075 , 
        \edb_top_inst/n1077 , \edb_top_inst/n1079 , \edb_top_inst/n1081 , 
        \edb_top_inst/n1083 , \edb_top_inst/n1085 , \edb_top_inst/n1087 , 
        \edb_top_inst/n1089 , \edb_top_inst/n1091 , \edb_top_inst/n1093 , 
        \edb_top_inst/n1095 , \edb_top_inst/n1097 , \edb_top_inst/n1099 , 
        \edb_top_inst/n1101 , \edb_top_inst/n1103 , \edb_top_inst/n1105 , 
        \edb_top_inst/n1107 , \edb_top_inst/n1109 , \edb_top_inst/n1111 , 
        \edb_top_inst/n1113 , \edb_top_inst/n1126 , \edb_top_inst/n1128 , 
        \edb_top_inst/n1130 , \edb_top_inst/n1132 , \edb_top_inst/n1134 , 
        \edb_top_inst/n1136 , \edb_top_inst/n1138 , \edb_top_inst/n1143 , 
        \edb_top_inst/n1145 , \edb_top_inst/n1147 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39] , 
        \edb_top_inst/n2758 , \edb_top_inst/n67 , \edb_top_inst/n1112 , 
        \edb_top_inst/n1110 , \edb_top_inst/n1108 , \edb_top_inst/n1106 , 
        \edb_top_inst/n1104 , \edb_top_inst/n1102 , \edb_top_inst/n1100 , 
        \edb_top_inst/n1098 , \edb_top_inst/n1096 , \edb_top_inst/n1094 , 
        \edb_top_inst/n1092 , \edb_top_inst/n1090 , \edb_top_inst/n1088 , 
        \edb_top_inst/n1086 , \edb_top_inst/n1084 , \edb_top_inst/n1082 , 
        \edb_top_inst/n1146 , \edb_top_inst/n1080 , \edb_top_inst/n1144 , 
        \edb_top_inst/n1078 , \edb_top_inst/n1142 , \edb_top_inst/n1076 , 
        \edb_top_inst/n1137 , \edb_top_inst/n1074 , \edb_top_inst/n1135 , 
        \edb_top_inst/n1072 , \edb_top_inst/n1133 , \edb_top_inst/n1070 , 
        \edb_top_inst/n1131 , \edb_top_inst/n1068 , \edb_top_inst/n1129 , 
        \edb_top_inst/n1066 , \edb_top_inst/n1127 , \edb_top_inst/n1064 , 
        \edb_top_inst/n1125 , \edb_top_inst/n1062 , \edb_top_inst/n1123 , 
        \edb_top_inst/n69 , \edb_top_inst/n1051 , \edb_top_inst/n1049 , 
        \edb_top_inst/n1047 , \edb_top_inst/n1046 , n9476, n9675, \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_1_q , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_0_q , n9759, 
        n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, 
        n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, 
        n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, 
        n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, 
        n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, 
        n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, 
        n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, 
        n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, 
        n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, 
        n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, 
        n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, 
        n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, 
        n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, 
        n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, 
        n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, 
        n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, 
        n9888, n9889, n9892, n9893, n9894, n9895, n9896, n9897, 
        n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, 
        n9906, n9913, n9914, n9915, n9916, n9917, n9918, n9919, 
        n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, 
        n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, 
        n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, 
        n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, 
        n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, 
        n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, 
        n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, 
        n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, 
        n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, 
        n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, 
        n10000, n10001, n10002, n10003, n10004, n10005, n10006, 
        n10007, n10008, n10009, n10010, n10011, n10012, n10013, 
        n10014, n10015, n10016, n10017, n10018, n10019, n10020, 
        n10021, n10022, n10023, n10024, n10025, n10026, n10027, 
        n10028, n10029, n10030, n10031, n10032, n10033, n10034, 
        n10035, n10036, n10037, n10038, n10039, n10040, n10041, 
        n10042, n10043, n10044, n10045, n10046, n10047, n10048, 
        n10049, n10050, n10051, n10052, n10053, n10054, n10055, 
        n10056, n10057, n10058, n10059, n10060, n10061, n10062, 
        n10063, n10064, n10065, n10066, n10067, n10068, n10069, 
        n10070, n10071, n10072, n10073, n10074, n10075, n10076, 
        n10077, n10078, n10079, n10080, n10081, n10082, n10083, 
        n10084, n10085, n10086, n10087, n10088, n10089, n10090, 
        n10091, n10092, n10093, n10094, n10095, n10096, n10097, 
        n10098, n10099, n10100, n10101, n10102, n10103, n10104, 
        n10105, n10106, n10107, n10108, n10109, n10110, n10111, 
        n10112, n10113, n10114, n10115, n10116, n10117, n10118, 
        n10119, n10120, n10121, n10122, n10123, n10124, n10125, 
        n10126, n10127, n10128, n10129, n10130, n10131, n10132, 
        n10133, n10134, n10135;
    
    assign MipiDphyRx1_RESET_N = MipiDphyRx1_RST0_N /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[2] = MipiDphyRx1_STOPSTATE_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign MipiDphyRx1_TX_REQUEST_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TURN_REQUEST = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_FORCE_RX_MODE = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_TRIGGER_ESC[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_TRIGGER_ESC[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_TRIGGER_ESC[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_TRIGGER_ESC[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[7] = MipiDphyRx1_RX_CLK_ACTIVE_HS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[10] = MipiDphyRx1_RX_ACTIVE_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[24] = MipiDphyRx1_RX_VALID_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[25] = MipiDphyRx1_RX_VALID_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[0] = MipiDphyRx1_RX_SYNC_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[3] = MipiDphyRx1_RX_SKEW_CAL_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[4] = MipiDphyRx1_RX_DATA_HS_LAN0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign MipiDphyRx1_TX_LPDT_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_VALID_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_READY_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_ULPS_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[17] = MipiDphyRx1_WORD_CLKOUT_HS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[1] = MipiDphyRx1_RX_CLK_ESC_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign MipiDphyRx1_TX_CLK_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oLed[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign pll_inst1_RSTN = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign pll_ddr_RSTN = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[23] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[22] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[21] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[20] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[19] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[18] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[16] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[15] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[14] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[13] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[12] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[11] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[9] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[8] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign jtag_inst1_TDO = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign pll_inst2_RSTN = 1'b1 /* verific EFX_ATTRIBUTE_CELL_NAME=VCC */ ;
    assign MipiDphyRx1_TX_ULPS_EXIT = 1'b0 /* verific EFX_ATTRIBUTE_CELL_NAME=GND */ ;
    EFX_FF \la0_probe4~FF  (.D(MipiDphyRx1_RX_SKEW_CAL_HS_LAN0), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(la0_probe4)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(288)
    defparam \la0_probe4~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe4~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe4~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe4~FF .D_POLARITY = 1'b1;
    defparam \la0_probe4~FF .SR_SYNC = 1'b0;
    defparam \la0_probe4~FF .SR_VALUE = 1'b0;
    defparam \la0_probe4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe10~FF  (.D(oTestPort[10]), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(la0_probe10)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(285)
    defparam \la0_probe10~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe10~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe10~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe10~FF .D_POLARITY = 1'b1;
    defparam \la0_probe10~FF .SR_SYNC = 1'b0;
    defparam \la0_probe10~FF .SR_VALUE = 1'b0;
    defparam \la0_probe10~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MipiDphyRx1_RESET_N~FF  (.D(oLed[5]), .CE(1'b1), .CLK(iSCLK), 
           .SR(iPushSw[0]), .Q(MipiDphyRx1_RST0_N)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MTopTi180MIPI25GRxHDMIV101.v(267)
    defparam \MipiDphyRx1_RESET_N~FF .CLK_POLARITY = 1'b1;
    defparam \MipiDphyRx1_RESET_N~FF .CE_POLARITY = 1'b1;
    defparam \MipiDphyRx1_RESET_N~FF .SR_POLARITY = 1'b0;
    defparam \MipiDphyRx1_RESET_N~FF .D_POLARITY = 1'b1;
    defparam \MipiDphyRx1_RESET_N~FF .SR_SYNC = 1'b0;
    defparam \MipiDphyRx1_RESET_N~FF .SR_VALUE = 1'b0;
    defparam \MipiDphyRx1_RESET_N~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rFRST~FF  (.D(oLed[5]), .CE(1'b1), .CLK(iFCLK), .SR(iPushSw[0]), 
           .Q(rFRST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MTopTi180MIPI25GRxHDMIV101.v(285)
    defparam \rFRST~FF .CLK_POLARITY = 1'b1;
    defparam \rFRST~FF .CE_POLARITY = 1'b1;
    defparam \rFRST~FF .SR_POLARITY = 1'b0;
    defparam \rFRST~FF .D_POLARITY = 1'b0;
    defparam \rFRST~FF .SR_SYNC = 1'b0;
    defparam \rFRST~FF .SR_VALUE = 1'b1;
    defparam \rFRST~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rBRST~FF  (.D(oLed[5]), .CE(1'b1), .CLK(iBCLK), .SR(iPushSw[0]), 
           .Q(rBRST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MTopTi180MIPI25GRxHDMIV101.v(296)
    defparam \rBRST~FF .CLK_POLARITY = 1'b1;
    defparam \rBRST~FF .CE_POLARITY = 1'b1;
    defparam \rBRST~FF .SR_POLARITY = 1'b0;
    defparam \rBRST~FF .D_POLARITY = 1'b0;
    defparam \rBRST~FF .SR_SYNC = 1'b0;
    defparam \rBRST~FF .SR_VALUE = 1'b1;
    defparam \rBRST~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rVRST~FF  (.D(oLed[5]), .CE(1'b1), .CLK(iVCLK), .SR(iPushSw[0]), 
           .Q(rVRST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MTopTi180MIPI25GRxHDMIV101.v(307)
    defparam \rVRST~FF .CLK_POLARITY = 1'b1;
    defparam \rVRST~FF .CE_POLARITY = 1'b1;
    defparam \rVRST~FF .SR_POLARITY = 1'b0;
    defparam \rVRST~FF .D_POLARITY = 1'b0;
    defparam \rVRST~FF .SR_SYNC = 1'b0;
    defparam \rVRST~FF .SR_VALUE = 1'b1;
    defparam \rVRST~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rnVRST~FF  (.D(oLed[5]), .CE(1'b1), .CLK(iVCLK), .SR(iPushSw[0]), 
           .Q(rnVRST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MTopTi180MIPI25GRxHDMIV101.v(311)
    defparam \rnVRST~FF .CLK_POLARITY = 1'b1;
    defparam \rnVRST~FF .CE_POLARITY = 1'b1;
    defparam \rnVRST~FF .SR_POLARITY = 1'b0;
    defparam \rnVRST~FF .D_POLARITY = 1'b1;
    defparam \rnVRST~FF .SR_SYNC = 1'b0;
    defparam \rnVRST~FF .SR_VALUE = 1'b0;
    defparam \rnVRST~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oLed[2]~FF  (.D(1'b1), .CE(wCdcFifoFull), .CLK(iSCLK), .SR(rSRST), 
           .Q(oLed[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MTopTi180MIPI25GRxHDMIV101.v(588)
    defparam \oLed[2]~FF .CLK_POLARITY = 1'b1;
    defparam \oLed[2]~FF .CE_POLARITY = 1'b1;
    defparam \oLed[2]~FF .SR_POLARITY = 1'b1;
    defparam \oLed[2]~FF .D_POLARITY = 1'b1;
    defparam \oLed[2]~FF .SR_SYNC = 1'b1;
    defparam \oLed[2]~FF .SR_VALUE = 1'b0;
    defparam \oLed[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe2~FF  (.D(MipiDphyRx1_STOPSTATE_LAN0), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(la0_probe2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(282)
    defparam \la0_probe2~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe2~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe2~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe2~FF .D_POLARITY = 1'b1;
    defparam \la0_probe2~FF .SR_SYNC = 1'b0;
    defparam \la0_probe2~FF .SR_VALUE = 1'b0;
    defparam \la0_probe2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe11~FF  (.D(oTestPort[24]), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(la0_probe11)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(279)
    defparam \la0_probe11~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe11~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe11~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe11~FF .D_POLARITY = 1'b1;
    defparam \la0_probe11~FF .SR_SYNC = 1'b0;
    defparam \la0_probe11~FF .SR_VALUE = 1'b0;
    defparam \la0_probe11~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[0]~FF  (.D(\MCsiRxController/n279 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[0]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[0]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[0]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[0]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[0]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[0]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[0]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[0]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(276)
    defparam \la0_probe9[0]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[0]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[0]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[0]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[0]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[0]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/n630 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/n632 ), 
           .Q(\MCsiRxController/MCsi2Decoder/rHsSt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(212)
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe3[0]~FF  (.D(oTestPort[0]), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe3[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe3[0]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe3[0]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe3[0]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe3[0]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe3[0]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe3[0]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe3[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF  (.D(\MCsiRxController/MCsi2Decoder/n7 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rSRST_2~FF  (.D(oLed[5]), .CE(1'b1), .CLK(iSCLK), .SR(iPushSw[0]), 
           .Q(rSRST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MTopTi180MIPI25GRxHDMIV101.v(263)
    defparam \rSRST_2~FF .CLK_POLARITY = 1'b1;
    defparam \rSRST_2~FF .CE_POLARITY = 1'b1;
    defparam \rSRST_2~FF .SR_POLARITY = 1'b0;
    defparam \rSRST_2~FF .D_POLARITY = 1'b0;
    defparam \rSRST_2~FF .SR_SYNC = 1'b0;
    defparam \rSRST_2~FF .SR_VALUE = 1'b1;
    defparam \rSRST_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe5~FF  (.D(MipiDphyRx1_ERR_SOT_HS_LAN0), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(la0_probe5)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(291)
    defparam \la0_probe5~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe5~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe5~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe5~FF .D_POLARITY = 1'b1;
    defparam \la0_probe5~FF .SR_SYNC = 1'b0;
    defparam \la0_probe5~FF .SR_VALUE = 1'b0;
    defparam \la0_probe5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe7~FF  (.D(MipiDphyRx1_RX_ERR_SYNC_ESC), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(la0_probe7)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(294)
    defparam \la0_probe7~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe7~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe7~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe7~FF .D_POLARITY = 1'b1;
    defparam \la0_probe7~FF .SR_SYNC = 1'b0;
    defparam \la0_probe7~FF .SR_VALUE = 1'b0;
    defparam \la0_probe7~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe0~FF  (.D(la0_probe0), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(la0_probe0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(264)
    defparam \la0_probe0~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe0~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe0~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe0~FF .D_POLARITY = 1'b0;
    defparam \la0_probe0~FF .SR_SYNC = 1'b0;
    defparam \la0_probe0~FF .SR_VALUE = 1'b0;
    defparam \la0_probe0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRVd ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(115)
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsValid~FF  (.D(\~MCsiRxController/MCsi2Decoder/reduce_nor_75/n1 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsValid )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsValid~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsValid~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsValid~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsValid~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/wHsValid~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsValid~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsValid~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/n603 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/n96 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\MCsiRxController/MCsi2Decoder/rHsSt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(212)
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/n606 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/n632 ), 
           .Q(\MCsiRxController/MCsi2Decoder/rHsSt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(212)
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[7]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[7]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe9[7]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[7]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[7]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[7]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[7]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[7]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[6]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[6]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe9[6]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[6]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[6]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[6]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[6]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[6]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[5]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[5]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe9[5]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[5]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[5]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[5]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[5]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[5]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[4]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[4]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe9[4]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[4]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[4]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[4]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[4]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[4]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[3]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[3]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe9[3]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[3]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[3]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[3]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[3]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[3]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[2]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[2]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe9[2]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[2]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[2]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[2]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[2]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[2]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[1]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[1]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe9[1]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[1]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[1]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[1]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[1]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[1]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/equal_38/n19 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/wFtiEmp[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(112)
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .SR_VALUE = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF  (.D(n117), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF  (.D(n3799), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF  (.D(n3797), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF  (.D(n3795), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF  (.D(n3793), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF  (.D(n3791), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF  (.D(n3789), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF  (.D(n3787), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF  (.D(n3786), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n233 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n238 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n243 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n248 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n253 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n258 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n263 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n268 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n273 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF  (.D(n120), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF  (.D(n169), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF  (.D(n3763), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF  (.D(n3761), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF  (.D(n3759), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF  (.D(n3757), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF  (.D(n3755), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF  (.D(n3753), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF  (.D(n3752), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[2] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[3] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[4] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[5] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[6] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[7] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[8]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[8] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[9]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[9] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[10]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[10] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[11]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[11] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[12]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[12] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[13]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[13] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[13]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[14]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[14] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[14]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[15]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[15] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/wHsPixel[15]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[9] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_62/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[1]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[1]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[1]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[10] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_62/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[2]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[2]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[2]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[11] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_62/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[3]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[3]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[3]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[12] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_62/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[4]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[4]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[4]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[13] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_62/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[5]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[5]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[5]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[14] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_62/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[6]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[6]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[6]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[15] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_62/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[7]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[7]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[7]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[8]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_59/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[8]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[8]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[8]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[8]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[9]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[1] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_59/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[9]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[9]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[9]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[9]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[10]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[2] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_59/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[10]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[10]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[10]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[10]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[11]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[3] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_59/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[11]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[11]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[11]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[11]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[12]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[4] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_59/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[12]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[12]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[12]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[12]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[12]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[13]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[5] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_59/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[13]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[13]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[13]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[13]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[13]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[14]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[6] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_59/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[14]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[14]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[14]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[14]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[14]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[15]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[7] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_59/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsWordCnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[15]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[15]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[15]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[15]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[15]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsDatatype[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[2] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_62/n5 ), .CLK(iSCLK), 
           .SR(rSRST), .Q(\wHsDatatype[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsDatatype[2]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsDatatype[2]~FF .CE_POLARITY = 1'b0;
    defparam \wHsDatatype[2]~FF .SR_POLARITY = 1'b1;
    defparam \wHsDatatype[2]~FF .D_POLARITY = 1'b1;
    defparam \wHsDatatype[2]~FF .SR_SYNC = 1'b1;
    defparam \wHsDatatype[2]~FF .SR_VALUE = 1'b0;
    defparam \wHsDatatype[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsDatatype[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[3] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_62/n5 ), .CLK(iSCLK), 
           .SR(rSRST), .Q(\wHsDatatype[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsDatatype[3]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsDatatype[3]~FF .CE_POLARITY = 1'b0;
    defparam \wHsDatatype[3]~FF .SR_POLARITY = 1'b1;
    defparam \wHsDatatype[3]~FF .D_POLARITY = 1'b1;
    defparam \wHsDatatype[3]~FF .SR_SYNC = 1'b1;
    defparam \wHsDatatype[3]~FF .SR_VALUE = 1'b0;
    defparam \wHsDatatype[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsDatatype[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[4] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_62/n5 ), .CLK(iSCLK), 
           .SR(rSRST), .Q(\wHsDatatype[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsDatatype[4]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsDatatype[4]~FF .CE_POLARITY = 1'b0;
    defparam \wHsDatatype[4]~FF .SR_POLARITY = 1'b1;
    defparam \wHsDatatype[4]~FF .D_POLARITY = 1'b1;
    defparam \wHsDatatype[4]~FF .SR_SYNC = 1'b1;
    defparam \wHsDatatype[4]~FF .SR_VALUE = 1'b0;
    defparam \wHsDatatype[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsDatatype[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[5] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_62/n5 ), .CLK(iSCLK), 
           .SR(rSRST), .Q(\wHsDatatype[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \wHsDatatype[5]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsDatatype[5]~FF .CE_POLARITY = 1'b0;
    defparam \wHsDatatype[5]~FF .SR_POLARITY = 1'b1;
    defparam \wHsDatatype[5]~FF .D_POLARITY = 1'b1;
    defparam \wHsDatatype[5]~FF .SR_SYNC = 1'b1;
    defparam \wHsDatatype[5]~FF .SR_VALUE = 1'b0;
    defparam \wHsDatatype[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF  (.D(n124), 
           .CE(\MCsiRxController/MCsi2Decoder/n603 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF  (.D(n3784), 
           .CE(\MCsiRxController/MCsi2Decoder/n603 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF  (.D(n3782), 
           .CE(\MCsiRxController/MCsi2Decoder/n603 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF  (.D(n3780), 
           .CE(\MCsiRxController/MCsi2Decoder/n603 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF  (.D(n3778), 
           .CE(\MCsiRxController/MCsi2Decoder/n603 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF  (.D(n3776), 
           .CE(\MCsiRxController/MCsi2Decoder/n603 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF  (.D(n3774), 
           .CE(\MCsiRxController/MCsi2Decoder/n603 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF  (.D(n3772), 
           .CE(\MCsiRxController/MCsi2Decoder/n603 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF  (.D(n3770), 
           .CE(\MCsiRxController/MCsi2Decoder/n603 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF  (.D(n3768), 
           .CE(\MCsiRxController/MCsi2Decoder/n603 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF  (.D(n3766), 
           .CE(\MCsiRxController/MCsi2Decoder/n603 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF  (.D(n3765), 
           .CE(\MCsiRxController/MCsi2Decoder/n603 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(273)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[0]~FF  (.D(oTestPort[4]), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe8[0]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[0]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[0]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[0]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[0]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[0]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[1]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[1]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe8[1]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[1]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[1]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[1]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[1]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[1]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[2]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[2]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe8[2]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[2]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[2]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[2]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[2]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[2]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[3]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[3]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe8[3]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[3]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[3]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[3]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[3]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[3]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[4]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[4]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe8[4]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[4]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[4]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[4]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[4]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[4]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[5]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[5]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe8[5]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[5]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[5]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[5]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[5]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[5]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[6]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[6]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe8[6]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[6]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[6]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[6]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[6]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[6]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[7]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[7]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(126)
    defparam \la0_probe8[7]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[7]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[7]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[7]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[7]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[7]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wCdcFifoFull_2~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/qFullAllmost ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(wCdcFifoFull)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(85)
    defparam \wCdcFifoFull_2~FF .CLK_POLARITY = 1'b1;
    defparam \wCdcFifoFull_2~FF .CE_POLARITY = 1'b1;
    defparam \wCdcFifoFull_2~FF .SR_POLARITY = 1'b0;
    defparam \wCdcFifoFull_2~FF .D_POLARITY = 1'b1;
    defparam \wCdcFifoFull_2~FF .SR_SYNC = 1'b0;
    defparam \wCdcFifoFull_2~FF .SR_VALUE = 1'b0;
    defparam \wCdcFifoFull_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wVideoVd~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/qRVD ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(wVideoVd)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(91)
    defparam \wVideoVd~FF .CLK_POLARITY = 1'b1;
    defparam \wVideoVd~FF .CE_POLARITY = 1'b1;
    defparam \wVideoVd~FF .SR_POLARITY = 1'b0;
    defparam \wVideoVd~FF .D_POLARITY = 1'b1;
    defparam \wVideoVd~FF .SR_SYNC = 1'b0;
    defparam \wVideoVd~FF .SR_VALUE = 1'b0;
    defparam \wVideoVd~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wFtiEmp[0]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/equal_75/n17 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/wFtiEmp[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(88)
    defparam \MCsiRxController/wFtiEmp[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wFtiEmp[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wFtiEmp[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/wFtiEmp[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/wFtiEmp[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/wFtiEmp[0]~FF .SR_VALUE = 1'b1;
    defparam \MCsiRxController/wFtiEmp[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF  (.D(n189), .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF  (.D(n210), .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF  (.D(n3750), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF  (.D(n3748), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF  (.D(n3746), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF  (.D(n3744), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF  (.D(n3742), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF  (.D(n3741), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n436 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n441 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n446 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n451 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n456 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n461 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n466 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n471 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[1]~FF  (.D(\MCsiRxController/n278 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[1]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[1]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[1]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[1]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[1]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[1]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[2]~FF  (.D(\MCsiRxController/n277 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[2]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[2]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[2]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[2]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[2]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[2]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[3]~FF  (.D(\MCsiRxController/n276 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[3]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[3]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[3]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[3]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[3]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[3]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[4]~FF  (.D(\MCsiRxController/n275 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[4]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[4]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[4]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[4]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[4]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[4]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[5]~FF  (.D(\MCsiRxController/n274 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[5]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[5]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[5]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[5]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[5]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[5]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[6]~FF  (.D(\MCsiRxController/n273 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[6]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[6]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[6]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[6]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[6]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[6]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[7]~FF  (.D(\MCsiRxController/n272 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[7]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[7]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[7]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[7]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[7]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[7]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[8]~FF  (.D(\MCsiRxController/n271 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[8]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[8]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[8]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[8]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[8]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[8]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[9]~FF  (.D(\MCsiRxController/n270 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[9]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[9]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[9]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[9]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[9]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[9]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[10]~FF  (.D(\MCsiRxController/n269 ), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[10]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[10]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[10]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[10]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[10]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[10]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[11]~FF  (.D(\MCsiRxController/n268 ), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[11]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[11]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[11]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[11]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[11]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[11]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[12]~FF  (.D(\MCsiRxController/n267 ), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[12]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[12]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[12]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[12]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[12]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[12]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[13]~FF  (.D(\MCsiRxController/n266 ), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[13]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[13]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[13]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[13]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[13]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[13]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[14]~FF  (.D(\MCsiRxController/n265 ), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[14]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[14]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[14]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[14]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[14]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[14]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[15]~FF  (.D(\MCsiRxController/n264 ), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe6[15]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[15]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[15]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[15]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[15]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[15]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe3[1]~FF  (.D(MipiDphyRx1_RX_SYNC_HS_LAN1), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe3[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(270)
    defparam \la0_probe3[1]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe3[1]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe3[1]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe3[1]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe3[1]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe3[1]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe3[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[0]~FF  (.D(\MVideoPostProcess/rVtgRstCnt[0] ), 
           .CE(\MVideoPostProcess/qVtgRstCntCke ), .CLK(iVCLK), .SR(rVRST), 
           .Q(\MVideoPostProcess/rVtgRstCnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRST[0]~FF  (.D(\MVideoPostProcess/rVtgRstSel ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRST[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRST[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstSel_2~FF  (.D(1'b0), .CE(\MVideoPostProcess/equal_18/n21 ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstSel )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF  (.D(\~n1834 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n816 ), 
           .CE(\~ceg_net512 ), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n833 ), 
           .CE(\~ceg_net512 ), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_last_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n268 ), 
           .CE(ceg_net995), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n277 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n242 ), 
           .CE(ceg_net1327), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15] ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1243 ), .CLK(iBCLK), 
           .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_2P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_clk_div_2P ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1243 ), .CLK(iBCLK), 
           .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_3P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n846 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n852 ), 
           .CE(ceg_net1087), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511SdaOe~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n847 ), 
           .CE(ceg_net1335), .CLK(iBCLK), .SR(rBRST), .Q(oAdv7511SdaOe)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \oAdv7511SdaOe~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511SdaOe~FF .CE_POLARITY = 1'b0;
    defparam \oAdv7511SdaOe~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511SdaOe~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511SdaOe~FF .SR_SYNC = 1'b0;
    defparam \oAdv7511SdaOe~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511SdaOe~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511SclOe~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n848 ), 
           .CE(ceg_net566), .CLK(iBCLK), .SR(rBRST), .Q(oAdv7511SclOe)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \oAdv7511SclOe~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511SclOe~FF .CE_POLARITY = 1'b0;
    defparam \oAdv7511SclOe~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511SclOe~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511SclOe~FF .SR_SYNC = 1'b0;
    defparam \oAdv7511SclOe~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511SclOe~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n870 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n879 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n829 ), 
           .CE(ceg_net1361), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/w_ack~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n899 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/w_ack )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n898 ), 
           .CE(ceg_net616), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n845 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n844 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n843 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n842 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n841 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n840 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n839 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n851 ), 
           .CE(ceg_net1087), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n850 ), 
           .CE(ceg_net1087), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n869 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n868 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n867 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n866 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n865 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n864 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n863 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n878 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n877 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n876 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n875 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n874 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n873 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n872 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n828 ), 
           .CE(ceg_net1471), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n827 ), 
           .CE(ceg_net1480), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n826 ), 
           .CE(ceg_net1488), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
            .I1(1'b1), .CI(1'b0), .CO(n10139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4659)
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[0] ), 
            .I1(1'b1), .CI(1'b0), .CO(n10138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4673)
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__MVideoPostProcess/mVideoTimingGen/add_6/i4  (.I0(n9675), 
            .I1(1'b1), .CI(1'b0), .CO(n10137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \AUX_ADD_CI__MVideoPostProcess/mVideoTimingGen/add_6/i4 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__MVideoPostProcess/mVideoTimingGen/add_6/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__genblk1.genblk1[0].mPulseGenerator/add_8/i4  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_1_q ), 
            .I1(1'b1), .CI(1'b0), .CO(n10136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \AUX_ADD_CI__genblk1.genblk1[0].mPulseGenerator/add_8/i4 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__genblk1.genblk1[0].mPulseGenerator/add_8/i4 .I1_POLARITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF  (.D(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2 ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF  (.D(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1 ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n251 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n250 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n249 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n248 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n247 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n246 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n245 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n244 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n700 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n705 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n710 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n715 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n720 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n725 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n730 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n735 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n740 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n745 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n750 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n755 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n760 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n765 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n770 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n780 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n785 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n790 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n795 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n800 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n805 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n810 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n276 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n275 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n274 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n273 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n272 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n271 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n270 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
           .CE(ceg_net1327), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n131 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/qVde ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/rVde[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(120)
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rHpos[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511Hs~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rHSync[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(oAdv7511Hs)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \oAdv7511Hs~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511Hs~FF .CE_POLARITY = 1'b1;
    defparam \oAdv7511Hs~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511Hs~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511Hs~FF .SR_SYNC = 1'b1;
    defparam \oAdv7511Hs~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511Hs~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n130 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n129 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF  (.D(n3697), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF  (.D(n3695), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n126 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n125 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF  (.D(n3689), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF  (.D(n3687), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF  (.D(n3685), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n121 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF  (.D(n3682), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511Vs~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rVSync[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(oAdv7511Vs)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \oAdv7511Vs~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511Vs~FF .CE_POLARITY = 1'b1;
    defparam \oAdv7511Vs~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511Vs~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511Vs~FF .SR_SYNC = 1'b1;
    defparam \oAdv7511Vs~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511Vs~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rVde[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/rVde[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(120)
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF  (.D(\MVideoPostProcess/wVgaGenFDe ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/rVde[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(120)
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511De~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rVde[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(oAdv7511De)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(120)
    defparam \oAdv7511De~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511De~FF .CE_POLARITY = 1'b1;
    defparam \oAdv7511De~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511De~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511De~FF .SR_SYNC = 1'b1;
    defparam \oAdv7511De~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511De~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/wVgaGenFDe_2~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rVde[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/wVgaGenFDe )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(120)
    defparam \MVideoPostProcess/wVgaGenFDe_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/wVgaGenFDe_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF  (.D(n436), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF  (.D(n3718), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF  (.D(n3716), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF  (.D(n3714), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF  (.D(n3712), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF  (.D(n3710), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF  (.D(n3708), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF  (.D(n3706), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF  (.D(n3704), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF  (.D(n3702), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF  (.D(n3701), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wVideofull~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qFullAllmost ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(wVideofull)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(105)
    defparam \wVideofull~FF .CLK_POLARITY = 1'b1;
    defparam \wVideofull~FF .CE_POLARITY = 1'b1;
    defparam \wVideofull~FF .SR_POLARITY = 1'b0;
    defparam \wVideofull~FF .D_POLARITY = 1'b1;
    defparam \wVideofull~FF .SR_SYNC = 1'b0;
    defparam \wVideofull~FF .SR_VALUE = 1'b0;
    defparam \wVideofull~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n495), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n3680), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3678), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3676), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3674), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3672), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3670), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3668), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3666), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3664), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3662), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3661), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF  (.D(\MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0 ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n478 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n483 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n488 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n493 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n498 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n503 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n508 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n513 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n518 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n523 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n528 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n533 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n560), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n532), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3659), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3657), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3655), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3653), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3651), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3649), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3647), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3645), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3643), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3642), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n604), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n577), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3640), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3638), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3636), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3634), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3632), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3630), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3628), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3626), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3624), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3623), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n648), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n621), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3621), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3619), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3617), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3615), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3613), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3611), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3609), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3607), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3605), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3604), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n692), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n665), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3602), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3600), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3598), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3596), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3594), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3592), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3590), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3588), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3586), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3585), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n736), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n709), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3583), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3581), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3579), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3577), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3575), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3573), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3571), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3569), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3567), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3566), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n780), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n753), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3564), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3562), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3560), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3558), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3556), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3554), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3552), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3550), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3548), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3547), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n824), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n797), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3545), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3543), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3541), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3539), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3537), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3535), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3533), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3531), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3529), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3528), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n868), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n841), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3526), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3524), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3522), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3520), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3518), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3516), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3514), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3512), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3510), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3509), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 LUT__13629 (.I0(\la0_probe6[0] ), .I1(oTestPort[24]), .O(\MCsiRxController/n279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13629.LUTMASK = 16'h4444;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n912), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n885), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3507), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3505), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3503), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3501), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3499), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3497), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3495), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3493), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3491), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3490), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n956), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n929), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3488), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3486), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3484), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3482), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3480), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3478), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3476), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3474), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3472), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3471), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n1000), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n973), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3469), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3467), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3465), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3463), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3461), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3459), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3457), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3455), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3453), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3452), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n1044), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n1017), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3450), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3448), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3446), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3444), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3442), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3440), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3438), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3436), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3434), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3433), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n1088), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n1061), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3431), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3429), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3427), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3425), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3423), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3421), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3419), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3417), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3415), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3414), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n1132), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n1105), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3412), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3410), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3408), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3406), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3404), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3402), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3400), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3398), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3396), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3395), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n1176), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n1149), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3393), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3391), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3389), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3387), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3385), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3383), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3381), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3379), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3377), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3376), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[1]~FF  (.D(n295), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[2]~FF  (.D(n331), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[3]~FF  (.D(n3739), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[4]~FF  (.D(n3737), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[5]~FF  (.D(n3735), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[6]~FF  (.D(n3733), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[7]~FF  (.D(n3731), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[8]~FF  (.D(n3729), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[9]~FF  (.D(n3727), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[10]~FF  (.D(n3726), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRST[1]~FF  (.D(\MVideoPostProcess/rVtgRST[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRST[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRST[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRST[2]_2~FF  (.D(\MVideoPostProcess/rVtgRST[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRST[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF  (.D(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] ), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .D_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oLed[0]~FF  (.D(oLed[0]), .CE(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), 
           .CLK(iFCLK), .SR(rFRST), .Q(oLed[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(71)
    defparam \oLed[0]~FF .CLK_POLARITY = 1'b1;
    defparam \oLed[0]~FF .CE_POLARITY = 1'b0;
    defparam \oLed[0]~FF .SR_POLARITY = 1'b1;
    defparam \oLed[0]~FF .D_POLARITY = 1'b0;
    defparam \oLed[0]~FF .SR_SYNC = 1'b1;
    defparam \oLed[0]~FF .SR_VALUE = 1'b0;
    defparam \oLed[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF  (.D(wVideoVd), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[0].mPulseGenerator/rSft[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF  (.D(n1219), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF  (.D(n1193), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF  (.D(n3374), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF  (.D(n3372), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF  (.D(n3370), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF  (.D(n3368), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF  (.D(n3366), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF  (.D(n3364), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF  (.D(n3362), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF  (.D(n3360), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF  (.D(n3358), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[12]~FF  (.D(n3357), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[12]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[12]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[12]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[12]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[12]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[12]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF  (.D(\genblk1.genblk1[0].mPulseGenerator/rSft[0] ), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[0].mPulseGenerator/rSft[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF  (.D(\genblk1.genblk1[0].mPulseGenerator/rSft[1] ), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[0].mPulseGenerator/rSft[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF  (.D(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[0] ), 
           .CE(\genblk1.genblk1[3].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] ), .Q(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .D_POLARITY = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oLed[3]~FF  (.D(oLed[3]), .CE(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] ), 
           .CLK(iFCLK), .SR(rFRST), .Q(oLed[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(71)
    defparam \oLed[3]~FF .CLK_POLARITY = 1'b1;
    defparam \oLed[3]~FF .CE_POLARITY = 1'b1;
    defparam \oLed[3]~FF .SR_POLARITY = 1'b1;
    defparam \oLed[3]~FF .D_POLARITY = 1'b0;
    defparam \oLed[3]~FF .SR_SYNC = 1'b1;
    defparam \oLed[3]~FF .SR_VALUE = 1'b0;
    defparam \oLed[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF  (.D(wCdcFifoFull), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[3].mPulseGenerator/rSft[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF  (.D(\genblk1.genblk1[3].mPulseGenerator/n50 ), 
           .CE(\genblk1.genblk1[3].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] ), .Q(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF  (.D(\genblk1.genblk1[3].mPulseGenerator/rSft[0] ), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[3].mPulseGenerator/rSft[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF  (.D(\genblk1.genblk1[3].mPulseGenerator/rSft[1] ), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[3].mPulseGenerator/rSft[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF  (.D(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[0] ), 
           .CE(\genblk1.genblk1[4].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] ), .Q(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .D_POLARITY = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oLed[4]~FF  (.D(oLed[4]), .CE(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] ), 
           .CLK(iFCLK), .SR(rFRST), .Q(oLed[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(71)
    defparam \oLed[4]~FF .CLK_POLARITY = 1'b1;
    defparam \oLed[4]~FF .CE_POLARITY = 1'b1;
    defparam \oLed[4]~FF .SR_POLARITY = 1'b1;
    defparam \oLed[4]~FF .D_POLARITY = 1'b0;
    defparam \oLed[4]~FF .SR_SYNC = 1'b1;
    defparam \oLed[4]~FF .SR_VALUE = 1'b0;
    defparam \oLed[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF  (.D(wVideofull), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[4].mPulseGenerator/rSft[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF  (.D(\genblk1.genblk1[4].mPulseGenerator/n50 ), 
           .CE(\genblk1.genblk1[4].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] ), .Q(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF  (.D(\genblk1.genblk1[4].mPulseGenerator/rSft[0] ), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[4].mPulseGenerator/rSft[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF  (.D(\genblk1.genblk1[4].mPulseGenerator/rSft[1] ), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[4].mPulseGenerator/rSft[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig~FF  (.D(\edb_top_inst/la0/n1340 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_run_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig_imdt~FF  (.D(\edb_top_inst/la0/n1341 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig_imdt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_stop_trig~FF  (.D(\edb_top_inst/la0/n1342 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_stop_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_stop_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[0]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[0]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_soft_reset_in~FF  (.D(\edb_top_inst/la0/n1965 ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_soft_reset_in )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3683)
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[0]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[0] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[0]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/opcode[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/opcode[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[0]~FF  (.D(\edb_top_inst/la0/n2189 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/bit_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[0]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[0] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[0]~FF  (.D(\edb_top_inst/la0/n2466 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[0]~FF  (.D(\edb_top_inst/la0/module_next_state[0] ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/module_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3794)
    defparam \edb_top_inst/la0/module_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn_p1~FF  (.D(1'b1), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_soft_reset_in ), .Q(\edb_top_inst/la0/la_resetn_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4104)
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn~FF  (.D(\edb_top_inst/la0/la_resetn_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_soft_reset_in ), 
           .Q(\edb_top_inst/la0/la_resetn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4104)
    defparam \edb_top_inst/la0/la_resetn~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF  (.D(la0_probe0), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF  (.D(la0_probe1), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF  (.D(la0_probe2), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF  (.D(\la0_probe3[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5294 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5492 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF  (.D(la0_probe4), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF  (.D(la0_probe5), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6947 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF  (.D(\la0_probe6[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF  (.D(la0_probe7), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n8741 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF  (.D(\la0_probe8[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF  (.D(\la0_probe9[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n10527 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF  (.D(la0_probe10), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n11368 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF  (.D(la0_probe11), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n12201 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[0]~FF  (.D(\edb_top_inst/edb_user_dr[64] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[0]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[32]~FF  (.D(\edb_top_inst/edb_user_dr[32] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[33]~FF  (.D(\edb_top_inst/edb_user_dr[33] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[34]~FF  (.D(\edb_top_inst/edb_user_dr[34] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[35]~FF  (.D(\edb_top_inst/edb_user_dr[35] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[36]~FF  (.D(\edb_top_inst/edb_user_dr[36] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[37]~FF  (.D(\edb_top_inst/edb_user_dr[37] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[38]~FF  (.D(\edb_top_inst/edb_user_dr[38] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[39]~FF  (.D(\edb_top_inst/edb_user_dr[39] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[40]~FF  (.D(\edb_top_inst/edb_user_dr[40] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[41]~FF  (.D(\edb_top_inst/edb_user_dr[41] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[42]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[43]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[44]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[45]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[46]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[47]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[48]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[49]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[50]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[51]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[52]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[53]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[54]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[55]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[56]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[57]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[58]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[59]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[60]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[61]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[62]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[63]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[1]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[2]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[3]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[4]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[5]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[6]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[7]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[8]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[9]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[10]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[11]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[12]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[13]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[14]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[15]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[16]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[1]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[2]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[3]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[4]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[1]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[1] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[2]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[2] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[3]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[3] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[4]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[4] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[5]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[5] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[6]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[6] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[7]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[7] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[8]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[8] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[9]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[9] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[10]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[10] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[11]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[11] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[12]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[12] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[13]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[13] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[14]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[14] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[15]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[15] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[16]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[16] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[17]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[17] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[18]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[18] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[19]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[19] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[20]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[20] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[21]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[21] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[22]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[22] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[23]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[23] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[24]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[24] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[25]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[25] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[26]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[26] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[1]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/opcode[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/opcode[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[2]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/opcode[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/opcode[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[3]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/opcode[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/opcode[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[1]~FF  (.D(\edb_top_inst/la0/n2188 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/bit_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[2]~FF  (.D(\edb_top_inst/la0/n2187 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/bit_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[3]~FF  (.D(\edb_top_inst/la0/n2186 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/bit_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[4]~FF  (.D(\edb_top_inst/la0/n2185 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/bit_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[5]~FF  (.D(\edb_top_inst/la0/n2184 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/bit_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[1]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[1] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[2]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[2] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[3]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[3] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[4]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[4] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[5]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[5] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[6]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[6] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[7]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[7] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[8]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[8] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[9]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[9] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[10]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[10] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[11]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[11] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[12]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[12] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[13]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[13] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[14]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[14] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[15]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[15] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[1]~FF  (.D(\edb_top_inst/la0/n2465 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[2]~FF  (.D(\edb_top_inst/la0/n2464 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[3]~FF  (.D(\edb_top_inst/la0/n2463 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[4]~FF  (.D(\edb_top_inst/la0/n2462 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[5]~FF  (.D(\edb_top_inst/la0/n2461 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[6]~FF  (.D(\edb_top_inst/la0/n2460 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[7]~FF  (.D(\edb_top_inst/la0/n2459 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[8]~FF  (.D(\edb_top_inst/la0/n2458 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[9]~FF  (.D(\edb_top_inst/la0/n2457 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[10]~FF  (.D(\edb_top_inst/la0/n2456 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[11]~FF  (.D(\edb_top_inst/la0/n2455 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[12]~FF  (.D(\edb_top_inst/la0/n2454 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[13]~FF  (.D(\edb_top_inst/la0/n2453 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[14]~FF  (.D(\edb_top_inst/la0/n2452 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[15]~FF  (.D(\edb_top_inst/la0/n2451 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[16]~FF  (.D(\edb_top_inst/la0/n2450 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[17]~FF  (.D(\edb_top_inst/la0/n2449 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[18]~FF  (.D(\edb_top_inst/la0/n2448 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[19]~FF  (.D(\edb_top_inst/la0/n2447 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[20]~FF  (.D(\edb_top_inst/la0/n2446 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[21]~FF  (.D(\edb_top_inst/la0/n2445 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[22]~FF  (.D(\edb_top_inst/la0/n2444 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[23]~FF  (.D(\edb_top_inst/la0/n2443 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[24]~FF  (.D(\edb_top_inst/la0/n2442 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[25]~FF  (.D(\edb_top_inst/la0/n2441 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[26]~FF  (.D(\edb_top_inst/la0/n2440 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[27]~FF  (.D(\edb_top_inst/la0/n2439 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[28]~FF  (.D(\edb_top_inst/la0/n2438 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[29]~FF  (.D(\edb_top_inst/la0/n2437 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[30]~FF  (.D(\edb_top_inst/la0/n2436 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[31]~FF  (.D(\edb_top_inst/la0/n2435 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[32]~FF  (.D(\edb_top_inst/la0/n2434 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[33]~FF  (.D(\edb_top_inst/la0/n2433 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[34]~FF  (.D(\edb_top_inst/la0/n2432 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[35]~FF  (.D(\edb_top_inst/la0/n2431 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[36]~FF  (.D(\edb_top_inst/la0/n2430 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[37]~FF  (.D(\edb_top_inst/la0/n2429 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[38]~FF  (.D(\edb_top_inst/la0/n2428 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[39]~FF  (.D(\edb_top_inst/la0/n2427 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[40]~FF  (.D(\edb_top_inst/la0/n2426 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[41]~FF  (.D(\edb_top_inst/la0/n2425 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[42]~FF  (.D(\edb_top_inst/la0/n2424 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[43]~FF  (.D(\edb_top_inst/la0/n2423 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[44]~FF  (.D(\edb_top_inst/la0/n2422 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[45]~FF  (.D(\edb_top_inst/la0/n2421 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[46]~FF  (.D(\edb_top_inst/la0/n2420 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[47]~FF  (.D(\edb_top_inst/la0/n2419 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[48]~FF  (.D(\edb_top_inst/la0/n2418 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[49]~FF  (.D(\edb_top_inst/la0/n2417 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[50]~FF  (.D(\edb_top_inst/la0/n2416 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[51]~FF  (.D(\edb_top_inst/la0/n2415 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[52]~FF  (.D(\edb_top_inst/la0/n2414 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[53]~FF  (.D(\edb_top_inst/la0/n2413 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[54]~FF  (.D(\edb_top_inst/la0/n2412 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[55]~FF  (.D(\edb_top_inst/la0/n2411 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[56]~FF  (.D(\edb_top_inst/la0/n2410 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[57]~FF  (.D(\edb_top_inst/la0/n2409 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[58]~FF  (.D(\edb_top_inst/la0/n2408 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[59]~FF  (.D(\edb_top_inst/la0/n2407 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[60]~FF  (.D(\edb_top_inst/la0/n2406 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[61]~FF  (.D(\edb_top_inst/la0/n2405 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[62]~FF  (.D(\edb_top_inst/la0/n2404 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[63]~FF  (.D(\edb_top_inst/la0/n2403 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[1]~FF  (.D(\edb_top_inst/la0/module_next_state[1] ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/module_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3794)
    defparam \edb_top_inst/la0/module_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[2]~FF  (.D(\edb_top_inst/la0/module_next_state[2] ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/module_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3794)
    defparam \edb_top_inst/la0/module_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[3]~FF  (.D(\edb_top_inst/la0/module_next_state[3] ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/module_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3794)
    defparam \edb_top_inst/la0/module_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[0]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n150 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[1]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n149 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[2]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n148 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[3]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n147 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[4]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n146 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[5]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n145 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[6]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n144 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[7]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n143 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[8]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n142 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[9]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n141 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[10]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n140 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[11]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n139 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[12]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n138 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[13]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n137 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[14]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n136 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[15]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n135 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[16]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n134 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[17]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n133 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[18]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n132 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[19]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n131 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[20]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n130 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[21]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n129 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[22]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n128 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[23]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n127 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[24]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n126 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[25]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n125 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[26]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n124 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[27]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n123 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[28]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n122 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[29]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n121 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[30]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n120 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[31]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n119 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n2766 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n2766 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n2766 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF  (.D(1'b1), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5522)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n3599 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n3599 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n3599 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n4432 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n4432 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n4432 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF  (.D(\la0_probe3[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5279 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5279 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n5279 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5294 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5492 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n10 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/equal_9/n3 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n26 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n9 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6114 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6114 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6114 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6947 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6947 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF  (.D(\la0_probe6[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF  (.D(\la0_probe6[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF  (.D(\la0_probe6[3] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF  (.D(\la0_probe6[4] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF  (.D(\la0_probe6[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF  (.D(\la0_probe6[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF  (.D(\la0_probe6[7] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF  (.D(\la0_probe6[8] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF  (.D(\la0_probe6[9] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF  (.D(\la0_probe6[10] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF  (.D(\la0_probe6[11] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF  (.D(\la0_probe6[12] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF  (.D(\la0_probe6[13] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF  (.D(\la0_probe6[14] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF  (.D(\la0_probe6[15] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n7892 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n7892 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n7892 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n72 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n38 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n73 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/equal_9/n31 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n82 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n71 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n70 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n69 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n68 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n67 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n66 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n65 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n64 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n63 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n62 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n61 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n60 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n59 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n58 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n57 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n37 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n36 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n35 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n34 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n33 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n32 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n31 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n30 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n29 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n28 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n27 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n26 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n25 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n24 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n8741 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n8741 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF  (.D(\la0_probe8[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF  (.D(\la0_probe8[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF  (.D(\la0_probe8[3] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF  (.D(\la0_probe8[4] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF  (.D(\la0_probe8[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF  (.D(\la0_probe8[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF  (.D(\la0_probe8[7] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n9630 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n9630 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n9630 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF  (.D(\la0_probe9[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF  (.D(\la0_probe9[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF  (.D(\la0_probe9[3] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF  (.D(\la0_probe9[4] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF  (.D(\la0_probe9[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF  (.D(\la0_probe9[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF  (.D(\la0_probe9[7] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/equal_9/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n38 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n37 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n36 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n35 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n34 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n33 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n21 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n20 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n19 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n10527 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n10527 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/equal_9/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n38 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n37 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n36 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n35 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n34 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n33 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n21 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n19 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n11368 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n11368 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n12201 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n12201 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/tu_trigger~FF  (.D(\edb_top_inst/la0/trigger_tu/n89 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/tu_trigger )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5764)
    defparam \edb_top_inst/la0/tu_trigger~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[40]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[41]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[2]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[5]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[6]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[23]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[23] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[40]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[40] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[41]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[41] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5250)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5050)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF  (.D(\edb_top_inst/la0/la_run_trig_imdt ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5050)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5050)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/str_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5271)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5286)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5286)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5286)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5296)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5309)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5309)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5309)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_fsm_state[0] ), 
           .CE(\edb_top_inst/ceg_net351 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5433)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1300 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/n17781 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5250)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5250)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5250)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF  (.D(\edb_top_inst/la0/la_run_trig ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5050)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/biu_ready~FF  (.D(\edb_top_inst/la0/la_biu_inst/n382 ), 
           .CE(\edb_top_inst/ceg_net348 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/biu_ready )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5321)
    defparam \edb_top_inst/la0/biu_ready~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF  (.D(\edb_top_inst/la0/address_counter[15] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF  (.D(\edb_top_inst/la0/address_counter[16] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF  (.D(\edb_top_inst/la0/address_counter[17] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF  (.D(\edb_top_inst/la0/address_counter[18] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF  (.D(\edb_top_inst/la0/address_counter[19] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF  (.D(\edb_top_inst/la0/address_counter[20] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF  (.D(\edb_top_inst/la0/address_counter[21] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF  (.D(\edb_top_inst/la0/address_counter[22] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF  (.D(\edb_top_inst/la0/address_counter[23] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF  (.D(\edb_top_inst/la0/address_counter[24] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF  (.D(\edb_top_inst/la0/address_counter[25] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF  (.D(\edb_top_inst/la0/address_counter[26] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[1] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[2] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[3] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[4] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[5] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[6] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[7] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[8] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[9] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[10] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[11] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[12]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[12] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[13]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[13] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[14]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[14] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[15]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[15] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[16]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[16] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[17]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[17] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[18]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[18] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[19]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[19] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[20]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[20] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[21]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[21] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[22]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[22] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[23]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[23] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[24]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[24] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[25]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[25] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[26]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[26] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[27]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[27] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[28]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[28] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[29]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[29] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[30]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[30] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[31]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[31] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[32]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[32] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[33]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[33] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[34]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[34] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[35]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[35] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[36]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[36] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[37]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[37] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[38]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[38] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[39]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[39] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[40]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[40] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[41]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[41] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[42]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[42] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_fsm_state[1] ), 
           .CE(\edb_top_inst/ceg_net351 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5433)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[0]~FF  (.D(\edb_top_inst/la0/la_sample_cnt[0] ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_push ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/n2053 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF  (.D(\edb_top_inst/n73 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF  (.D(\edb_top_inst/n1044 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF  (.D(\edb_top_inst/n1042 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF  (.D(\edb_top_inst/n1040 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF  (.D(\edb_top_inst/n1038 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF  (.D(\edb_top_inst/n1036 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF  (.D(\edb_top_inst/n1034 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF  (.D(\edb_top_inst/n1032 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF  (.D(\edb_top_inst/n1030 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF  (.D(\edb_top_inst/n1028 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF  (.D(\edb_top_inst/n1027 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF  (.D(\edb_top_inst/n693 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF  (.D(\edb_top_inst/n1025 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF  (.D(\edb_top_inst/n1023 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF  (.D(\edb_top_inst/n1021 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF  (.D(\edb_top_inst/n1019 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF  (.D(\edb_top_inst/n1017 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF  (.D(\edb_top_inst/n1015 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF  (.D(\edb_top_inst/n1013 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF  (.D(\edb_top_inst/n1011 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF  (.D(\edb_top_inst/n1008 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF  (.D(\edb_top_inst/n1005 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF  (.D(\edb_top_inst/n695 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF  (.D(\edb_top_inst/n856 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF  (.D(\edb_top_inst/n854 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF  (.D(\edb_top_inst/n852 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF  (.D(\edb_top_inst/n850 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF  (.D(\edb_top_inst/n848 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF  (.D(\edb_top_inst/n846 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF  (.D(\edb_top_inst/n844 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF  (.D(\edb_top_inst/n842 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF  (.D(\edb_top_inst/n840 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF  (.D(\edb_top_inst/n838 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[1]~FF  (.D(\edb_top_inst/n710 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[2]~FF  (.D(\edb_top_inst/n731 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[3]~FF  (.D(\edb_top_inst/n729 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[4]~FF  (.D(\edb_top_inst/n727 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[5]~FF  (.D(\edb_top_inst/n725 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[6]~FF  (.D(\edb_top_inst/n723 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[7]~FF  (.D(\edb_top_inst/n721 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[8]~FF  (.D(\edb_top_inst/n719 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[9]~FF  (.D(\edb_top_inst/n717 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[10]~FF  (.D(\edb_top_inst/n715 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[11]~FF  (.D(\edb_top_inst/n713 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[12]~FF  (.D(\edb_top_inst/n712 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[23] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[40] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[41] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[11] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[11] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF  (.D(\edb_top_inst/n711 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF  (.D(\edb_top_inst/n752 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF  (.D(\edb_top_inst/n750 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF  (.D(\edb_top_inst/n748 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF  (.D(\edb_top_inst/n746 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF  (.D(\edb_top_inst/n744 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF  (.D(\edb_top_inst/n742 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF  (.D(\edb_top_inst/n740 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF  (.D(\edb_top_inst/n738 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF  (.D(\edb_top_inst/n736 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF  (.D(\edb_top_inst/n734 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF  (.D(\edb_top_inst/n733 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[1]~FF  (.D(\edb_top_inst/edb_user_dr[65] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[2]~FF  (.D(\edb_top_inst/edb_user_dr[66] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[3]~FF  (.D(\edb_top_inst/edb_user_dr[67] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[4]~FF  (.D(\edb_top_inst/edb_user_dr[68] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[5]~FF  (.D(\edb_top_inst/edb_user_dr[69] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[6]~FF  (.D(\edb_top_inst/edb_user_dr[70] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[7]~FF  (.D(\edb_top_inst/edb_user_dr[71] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[8]~FF  (.D(\edb_top_inst/edb_user_dr[72] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[9]~FF  (.D(\edb_top_inst/edb_user_dr[73] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[10]~FF  (.D(\edb_top_inst/edb_user_dr[74] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[11]~FF  (.D(\edb_top_inst/edb_user_dr[75] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[12]~FF  (.D(\edb_top_inst/edb_user_dr[76] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[1]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[2]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[3]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[4]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[5]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[6]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[7]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[8]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[9]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[10]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[11]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[12]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[13]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[14]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[15]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[16]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(355)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[0]_2~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(355)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(355)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(355)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[1]_2~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[2]_2~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[3]_2~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[4]_2~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[5]_2~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[6]_2~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[7]_2~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[8]_2~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[9]_2~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[10]_2~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[11]_2~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[12]_2~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[13]_2~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[14]_2~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[15]_2~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[16]_2~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[17]_2~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[18]_2~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[19]_2~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[20]_2~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[21]_2~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[22]_2~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[23]_2~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[24]_2~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[25]_2~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[26]_2~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[27]_2~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[28]_2~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[29]_2~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[30]_2~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[31]_2~FF  (.D(\edb_top_inst/edb_user_dr[32] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[32]_2~FF  (.D(\edb_top_inst/edb_user_dr[33] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[33]_2~FF  (.D(\edb_top_inst/edb_user_dr[34] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[34]_2~FF  (.D(\edb_top_inst/edb_user_dr[35] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[35]_2~FF  (.D(\edb_top_inst/edb_user_dr[36] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[36]_2~FF  (.D(\edb_top_inst/edb_user_dr[37] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[37]_2~FF  (.D(\edb_top_inst/edb_user_dr[38] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[38]_2~FF  (.D(\edb_top_inst/edb_user_dr[39] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[39]_2~FF  (.D(\edb_top_inst/edb_user_dr[40] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[40]_2~FF  (.D(\edb_top_inst/edb_user_dr[41] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[41]_2~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[42]_2~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[43]_2~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[44]_2~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[45]_2~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[46]_2~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[47]_2~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[48]_2~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[49]_2~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[50]_2~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[51]_2~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[52]_2~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[53]_2~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[54]_2~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[55]_2~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[56]_2~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[57]_2~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[58]_2~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[59]_2~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[60]_2~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[61]_2~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[62]_2~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[63]_2~FF  (.D(\edb_top_inst/edb_user_dr[64] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[64]_2~FF  (.D(\edb_top_inst/edb_user_dr[65] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[65]_2~FF  (.D(\edb_top_inst/edb_user_dr[66] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[66]_2~FF  (.D(\edb_top_inst/edb_user_dr[67] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[67]_2~FF  (.D(\edb_top_inst/edb_user_dr[68] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[68]_2~FF  (.D(\edb_top_inst/edb_user_dr[69] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[69]_2~FF  (.D(\edb_top_inst/edb_user_dr[70] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[70]_2~FF  (.D(\edb_top_inst/edb_user_dr[71] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[71]_2~FF  (.D(\edb_top_inst/edb_user_dr[72] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[72]_2~FF  (.D(\edb_top_inst/edb_user_dr[73] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[73]_2~FF  (.D(\edb_top_inst/edb_user_dr[74] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[74]_2~FF  (.D(\edb_top_inst/edb_user_dr[75] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[75]_2~FF  (.D(\edb_top_inst/edb_user_dr[76] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[76]_2~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[77]_2~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[78]_2~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[79]_2~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[80]_2~FF  (.D(\edb_top_inst/edb_user_dr[81] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[81]_2~FF  (.D(jtag_inst2_TDI), .CE(\edb_top_inst/debug_hub_inst/n95 ), 
           .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i2  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
            .CI(1'b0), .O(n117), .CO(n118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i2  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0] ), 
            .CI(1'b0), .O(n120), .CO(n121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_48/i2  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] ), .CI(1'b0), 
            .O(n124), .CO(n125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(269)
    defparam \MCsiRxController/MCsi2Decoder/add_48/i2 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_48/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i3  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I1(1'b0), .CI(n121), .O(n169), .CO(n170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i2  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), .CI(1'b0), 
            .O(n189), .CO(n190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i2 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i3  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n190), .O(n210), .CO(n211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i3 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i2  (.I0(\MVideoPostProcess/rVtgRstCnt[1] ), 
            .I1(\MVideoPostProcess/rVtgRstCnt[0] ), .CI(1'b0), .O(n295), 
            .CO(n296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i3  (.I0(\MVideoPostProcess/rVtgRstCnt[2] ), 
            .I1(1'b0), .CI(n296), .O(n331), .CO(n332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i2  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[1] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[0] ), .CI(1'b0), 
            .O(n436), .CO(n437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i2  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[1] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[0] ), .CI(1'b0), 
            .O(n492), .CO(n493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n495), .CO(n496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n561), .O(n532), .CO(n533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n560), .CO(n561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n605), .O(n577), .CO(n578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n604), .CO(n605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n649), .O(n621), .CO(n622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n648), .CO(n649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n693), .O(n665), .CO(n666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n692), .CO(n693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n737), .O(n709), .CO(n710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n736), .CO(n737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n781), .O(n753), .CO(n754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n780), .CO(n781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n825), .O(n797), .CO(n798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n824), .CO(n825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n869), .O(n841), .CO(n842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n868), .CO(n869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n913), .O(n885), .CO(n886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n912), .CO(n913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n957), .O(n929), .CO(n930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n956), .CO(n957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n1001), .O(n973), .CO(n974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n1000), .CO(n1001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n1045), .O(n1017), .CO(n1018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n1044), .CO(n1045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n1089), .O(n1061), .CO(n1062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n1088), .CO(n1089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n1133), .O(n1105), .CO(n1106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n1132), .CO(n1133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n1177), .O(n1149), .CO(n1150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n1176), .CO(n1177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i3  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[2] ), 
            .I1(1'b0), .CI(n1220), .O(n1193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i3 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i2  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[1] ), 
            .I1(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] ), .CI(1'b0), 
            .O(n1219), .CO(n1220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i2 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i13  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[12] ), 
            .I1(1'b0), .CI(n3359), .O(n3357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i13 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i12  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[11] ), 
            .I1(1'b0), .CI(n3361), .O(n3358), .CO(n3359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i12 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i11  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[10] ), 
            .I1(1'b0), .CI(n3363), .O(n3360), .CO(n3361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i11 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i10  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[9] ), 
            .I1(1'b0), .CI(n3365), .O(n3362), .CO(n3363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i10 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i9  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[8] ), 
            .I1(1'b0), .CI(n3367), .O(n3364), .CO(n3365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i9 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i8  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[7] ), 
            .I1(1'b0), .CI(n3369), .O(n3366), .CO(n3367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i8 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i7  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[6] ), 
            .I1(1'b0), .CI(n3371), .O(n3368), .CO(n3369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i7 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i6  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[5] ), 
            .I1(1'b0), .CI(n3373), .O(n3370), .CO(n3371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i6 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i5  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[4] ), 
            .I1(1'b0), .CI(n3375), .O(n3372), .CO(n3373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i5 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i4  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[3] ), 
            .I1(1'b0), .CI(n10136), .O(n3374), .CO(n3375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i4 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3378), .O(n3376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3380), .O(n3377), .CO(n3378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3382), .O(n3379), .CO(n3380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3384), .O(n3381), .CO(n3382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3386), .O(n3383), .CO(n3384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3388), .O(n3385), .CO(n3386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3390), .O(n3387), .CO(n3388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3392), .O(n3389), .CO(n3390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3394), .O(n3391), .CO(n3392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n1150), .O(n3393), .CO(n3394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3397), .O(n3395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3399), .O(n3396), .CO(n3397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3401), .O(n3398), .CO(n3399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3403), .O(n3400), .CO(n3401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3405), .O(n3402), .CO(n3403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3407), .O(n3404), .CO(n3405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3409), .O(n3406), .CO(n3407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3411), .O(n3408), .CO(n3409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3413), .O(n3410), .CO(n3411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n1106), .O(n3412), .CO(n3413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3416), .O(n3414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3418), .O(n3415), .CO(n3416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3420), .O(n3417), .CO(n3418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3422), .O(n3419), .CO(n3420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3424), .O(n3421), .CO(n3422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3426), .O(n3423), .CO(n3424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3428), .O(n3425), .CO(n3426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3430), .O(n3427), .CO(n3428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3432), .O(n3429), .CO(n3430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n1062), .O(n3431), .CO(n3432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3435), .O(n3433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3437), .O(n3434), .CO(n3435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3439), .O(n3436), .CO(n3437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3441), .O(n3438), .CO(n3439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3443), .O(n3440), .CO(n3441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3445), .O(n3442), .CO(n3443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3447), .O(n3444), .CO(n3445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3449), .O(n3446), .CO(n3447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3451), .O(n3448), .CO(n3449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n1018), .O(n3450), .CO(n3451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3454), .O(n3452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3456), .O(n3453), .CO(n3454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3458), .O(n3455), .CO(n3456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3460), .O(n3457), .CO(n3458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3462), .O(n3459), .CO(n3460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3464), .O(n3461), .CO(n3462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3466), .O(n3463), .CO(n3464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3468), .O(n3465), .CO(n3466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3470), .O(n3467), .CO(n3468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n974), .O(n3469), .CO(n3470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3473), .O(n3471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3475), .O(n3472), .CO(n3473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3477), .O(n3474), .CO(n3475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3479), .O(n3476), .CO(n3477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3481), .O(n3478), .CO(n3479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3483), .O(n3480), .CO(n3481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3485), .O(n3482), .CO(n3483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3487), .O(n3484), .CO(n3485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3489), .O(n3486), .CO(n3487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n930), .O(n3488), .CO(n3489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3492), .O(n3490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3494), .O(n3491), .CO(n3492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3496), .O(n3493), .CO(n3494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3498), .O(n3495), .CO(n3496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3500), .O(n3497), .CO(n3498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3502), .O(n3499), .CO(n3500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3504), .O(n3501), .CO(n3502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3506), .O(n3503), .CO(n3504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3508), .O(n3505), .CO(n3506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n886), .O(n3507), .CO(n3508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3511), .O(n3509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3513), .O(n3510), .CO(n3511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3515), .O(n3512), .CO(n3513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3517), .O(n3514), .CO(n3515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3519), .O(n3516), .CO(n3517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3521), .O(n3518), .CO(n3519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3523), .O(n3520), .CO(n3521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3525), .O(n3522), .CO(n3523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3527), .O(n3524), .CO(n3525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n842), .O(n3526), .CO(n3527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3530), .O(n3528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3532), .O(n3529), .CO(n3530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3534), .O(n3531), .CO(n3532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3536), .O(n3533), .CO(n3534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3538), .O(n3535), .CO(n3536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3540), .O(n3537), .CO(n3538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3542), .O(n3539), .CO(n3540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3544), .O(n3541), .CO(n3542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3546), .O(n3543), .CO(n3544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n798), .O(n3545), .CO(n3546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3549), .O(n3547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3551), .O(n3548), .CO(n3549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3553), .O(n3550), .CO(n3551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3555), .O(n3552), .CO(n3553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3557), .O(n3554), .CO(n3555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3559), .O(n3556), .CO(n3557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3561), .O(n3558), .CO(n3559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3563), .O(n3560), .CO(n3561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3565), .O(n3562), .CO(n3563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n754), .O(n3564), .CO(n3565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3568), .O(n3566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3570), .O(n3567), .CO(n3568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3572), .O(n3569), .CO(n3570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3574), .O(n3571), .CO(n3572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3576), .O(n3573), .CO(n3574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3578), .O(n3575), .CO(n3576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3580), .O(n3577), .CO(n3578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3582), .O(n3579), .CO(n3580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3584), .O(n3581), .CO(n3582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n710), .O(n3583), .CO(n3584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3587), .O(n3585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3589), .O(n3586), .CO(n3587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3591), .O(n3588), .CO(n3589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3593), .O(n3590), .CO(n3591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3595), .O(n3592), .CO(n3593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3597), .O(n3594), .CO(n3595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3599), .O(n3596), .CO(n3597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3601), .O(n3598), .CO(n3599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3603), .O(n3600), .CO(n3601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n666), .O(n3602), .CO(n3603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3606), .O(n3604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3608), .O(n3605), .CO(n3606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3610), .O(n3607), .CO(n3608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3612), .O(n3609), .CO(n3610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3614), .O(n3611), .CO(n3612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3616), .O(n3613), .CO(n3614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3618), .O(n3615), .CO(n3616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3620), .O(n3617), .CO(n3618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3622), .O(n3619), .CO(n3620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n622), .O(n3621), .CO(n3622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3625), .O(n3623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3627), .O(n3624), .CO(n3625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3629), .O(n3626), .CO(n3627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3631), .O(n3628), .CO(n3629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3633), .O(n3630), .CO(n3631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3635), .O(n3632), .CO(n3633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3637), .O(n3634), .CO(n3635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3639), .O(n3636), .CO(n3637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3641), .O(n3638), .CO(n3639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n578), .O(n3640), .CO(n3641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3644), .O(n3642)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3646), .O(n3643), .CO(n3644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3648), .O(n3645), .CO(n3646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3650), .O(n3647), .CO(n3648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3652), .O(n3649), .CO(n3650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3654), .O(n3651), .CO(n3652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3656), .O(n3653), .CO(n3654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3658), .O(n3655), .CO(n3656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3660), .O(n3657), .CO(n3658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n533), .O(n3659), .CO(n3660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3663), .O(n3661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3665), .O(n3662), .CO(n3663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3667), .O(n3664), .CO(n3665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3669), .O(n3666), .CO(n3667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3671), .O(n3668), .CO(n3669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3673), .O(n3670), .CO(n3671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3675), .O(n3672), .CO(n3673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3677), .O(n3674), .CO(n3675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3679), .O(n3676), .CO(n3677)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n3681), .O(n3678), .CO(n3679)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n496), .O(n3680), .CO(n3681)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i12  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[11] ), 
            .I1(1'b0), .CI(n3684), .O(n3682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i11  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[10] ), 
            .I1(1'b0), .CI(n3686), .O(n3683), .CO(n3684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i10  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[9] ), 
            .I1(1'b0), .CI(n3688), .O(n3685), .CO(n3686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i9  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[8] ), 
            .I1(1'b0), .CI(n3690), .O(n3687), .CO(n3688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i8  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[7] ), 
            .I1(1'b0), .CI(n3692), .O(n3689), .CO(n3690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i7  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[6] ), 
            .I1(1'b0), .CI(n3694), .O(n3691), .CO(n3692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i6  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[5] ), 
            .I1(1'b0), .CI(n3696), .O(n3693), .CO(n3694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i5  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[4] ), 
            .I1(1'b0), .CI(n3698), .O(n3695), .CO(n3696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i4  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[3] ), 
            .I1(1'b0), .CI(n3700), .O(n3697), .CO(n3698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i3  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[2] ), 
            .I1(1'b0), .CI(n493), .O(n3699), .CO(n3700)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i12  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[11] ), 
            .I1(1'b0), .CI(n3703), .O(n3701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i11  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[10] ), 
            .I1(1'b0), .CI(n3705), .O(n3702), .CO(n3703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i10  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[9] ), 
            .I1(1'b0), .CI(n3707), .O(n3704), .CO(n3705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i9  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[8] ), 
            .I1(1'b0), .CI(n3709), .O(n3706), .CO(n3707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i8  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[7] ), 
            .I1(1'b0), .CI(n3711), .O(n3708), .CO(n3709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i7  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[6] ), 
            .I1(1'b0), .CI(n3713), .O(n3710), .CO(n3711)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i6  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[5] ), 
            .I1(1'b0), .CI(n3715), .O(n3712), .CO(n3713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i5  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[4] ), 
            .I1(1'b0), .CI(n3717), .O(n3714), .CO(n3715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i4  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[3] ), 
            .I1(1'b0), .CI(n10137), .O(n3716), .CO(n3717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i3  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[2] ), 
            .I1(1'b0), .CI(n437), .O(n3718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i11  (.I0(\MVideoPostProcess/rVtgRstCnt[10] ), 
            .I1(1'b0), .CI(n3728), .O(n3726)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i10  (.I0(\MVideoPostProcess/rVtgRstCnt[9] ), 
            .I1(1'b0), .CI(n3730), .O(n3727), .CO(n3728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i9  (.I0(\MVideoPostProcess/rVtgRstCnt[8] ), 
            .I1(1'b0), .CI(n3732), .O(n3729), .CO(n3730)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i8  (.I0(\MVideoPostProcess/rVtgRstCnt[7] ), 
            .I1(1'b0), .CI(n3734), .O(n3731), .CO(n3732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i7  (.I0(\MVideoPostProcess/rVtgRstCnt[6] ), 
            .I1(1'b0), .CI(n3736), .O(n3733), .CO(n3734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i6  (.I0(\MVideoPostProcess/rVtgRstCnt[5] ), 
            .I1(1'b0), .CI(n3738), .O(n3735), .CO(n3736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i5  (.I0(\MVideoPostProcess/rVtgRstCnt[4] ), 
            .I1(1'b0), .CI(n3740), .O(n3737), .CO(n3738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i4  (.I0(\MVideoPostProcess/rVtgRstCnt[3] ), 
            .I1(1'b0), .CI(n332), .O(n3739), .CO(n3740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i9  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3743), .O(n3741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i9 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i8  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3745), .O(n3742), .CO(n3743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i8 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i7  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3747), .O(n3744), .CO(n3745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i7 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i6  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3749), .O(n3746), .CO(n3747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i6 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i5  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3751), .O(n3748), .CO(n3749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i5 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i4  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n211), .O(n3750), .CO(n3751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i4 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i10  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9] ), 
            .I1(1'b0), .CI(n3754), .O(n3752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i9  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8] ), 
            .I1(1'b0), .CI(n3756), .O(n3753), .CO(n3754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i8  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7] ), 
            .I1(1'b0), .CI(n3758), .O(n3755), .CO(n3756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i7  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6] ), 
            .I1(1'b0), .CI(n3760), .O(n3757), .CO(n3758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i6  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5] ), 
            .I1(1'b0), .CI(n3762), .O(n3759), .CO(n3760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i5  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4] ), 
            .I1(1'b0), .CI(n3764), .O(n3761), .CO(n3762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i4  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3] ), 
            .I1(1'b0), .CI(n170), .O(n3763), .CO(n3764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_48/i13  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12] ), 
            .I1(1'b0), .CI(n3767), .O(n3765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(269)
    defparam \MCsiRxController/MCsi2Decoder/add_48/i13 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_48/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_48/i12  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] ), 
            .I1(1'b0), .CI(n3769), .O(n3766), .CO(n3767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(269)
    defparam \MCsiRxController/MCsi2Decoder/add_48/i12 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_48/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_48/i11  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] ), 
            .I1(1'b0), .CI(n3771), .O(n3768), .CO(n3769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(269)
    defparam \MCsiRxController/MCsi2Decoder/add_48/i11 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_48/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_48/i10  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9] ), 
            .I1(1'b0), .CI(n3773), .O(n3770), .CO(n3771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(269)
    defparam \MCsiRxController/MCsi2Decoder/add_48/i10 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_48/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_48/i9  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8] ), 
            .I1(1'b0), .CI(n3775), .O(n3772), .CO(n3773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(269)
    defparam \MCsiRxController/MCsi2Decoder/add_48/i9 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_48/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_48/i8  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7] ), 
            .I1(1'b0), .CI(n3777), .O(n3774), .CO(n3775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(269)
    defparam \MCsiRxController/MCsi2Decoder/add_48/i8 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_48/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_48/i7  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6] ), 
            .I1(1'b0), .CI(n3779), .O(n3776), .CO(n3777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(269)
    defparam \MCsiRxController/MCsi2Decoder/add_48/i7 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_48/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_48/i6  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5] ), 
            .I1(1'b0), .CI(n3781), .O(n3778), .CO(n3779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(269)
    defparam \MCsiRxController/MCsi2Decoder/add_48/i6 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_48/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_48/i5  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4] ), 
            .I1(1'b0), .CI(n3783), .O(n3780), .CO(n3781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(269)
    defparam \MCsiRxController/MCsi2Decoder/add_48/i5 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_48/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_48/i4  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3] ), 
            .I1(1'b0), .CI(n3785), .O(n3782), .CO(n3783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(269)
    defparam \MCsiRxController/MCsi2Decoder/add_48/i4 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_48/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_48/i3  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2] ), 
            .I1(1'b0), .CI(n125), .O(n3784), .CO(n3785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(269)
    defparam \MCsiRxController/MCsi2Decoder/add_48/i3 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_48/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i10  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] ), 
            .I1(1'b0), .CI(n3788), .O(n3786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i9  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] ), 
            .I1(1'b0), .CI(n3790), .O(n3787), .CO(n3788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i8  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
            .I1(1'b0), .CI(n3792), .O(n3789), .CO(n3790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i7  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] ), 
            .I1(1'b0), .CI(n3794), .O(n3791), .CO(n3792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i6  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
            .I1(1'b0), .CI(n3796), .O(n3793), .CO(n3794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i5  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] ), 
            .I1(1'b0), .CI(n3798), .O(n3795), .CO(n3796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i4  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] ), 
            .I1(1'b0), .CI(n3800), .O(n3797), .CO(n3798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i3  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I1(1'b0), .CI(n118), .O(n3799), .CO(n3800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i16  (.I0(\la0_probe6[15] ), .I1(1'b0), 
            .CI(n3803), .O(n3801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i16 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i15  (.I0(\la0_probe6[14] ), .I1(1'b0), 
            .CI(n3805), .O(n3802), .CO(n3803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i15 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i14  (.I0(\la0_probe6[13] ), .I1(1'b0), 
            .CI(n3807), .O(n3804), .CO(n3805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i14 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i13  (.I0(\la0_probe6[12] ), .I1(1'b0), 
            .CI(n3809), .O(n3806), .CO(n3807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i13 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i12  (.I0(\la0_probe6[11] ), .I1(1'b0), 
            .CI(n3811), .O(n3808), .CO(n3809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i12 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i11  (.I0(\la0_probe6[10] ), .I1(1'b0), 
            .CI(n3813), .O(n3810), .CO(n3811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i11 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i10  (.I0(\la0_probe6[9] ), .I1(1'b0), 
            .CI(n3815), .O(n3812), .CO(n3813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i10 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i9  (.I0(\la0_probe6[8] ), .I1(1'b0), 
            .CI(n3817), .O(n3814), .CO(n3815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i9 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i8  (.I0(\la0_probe6[7] ), .I1(1'b0), 
            .CI(n3819), .O(n3816), .CO(n3817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i8 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i7  (.I0(\la0_probe6[6] ), .I1(1'b0), 
            .CI(n3821), .O(n3818), .CO(n3819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i7 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i6  (.I0(\la0_probe6[5] ), .I1(1'b0), 
            .CI(n3823), .O(n3820), .CO(n3821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i6 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i5  (.I0(\la0_probe6[4] ), .I1(1'b0), 
            .CI(n3825), .O(n3822), .CO(n3823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i5 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i4  (.I0(\la0_probe6[3] ), .I1(1'b0), 
            .CI(n3827), .O(n3824), .CO(n3825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i4 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i3  (.I0(\la0_probe6[2] ), .I1(1'b0), 
            .CI(n3829), .O(n3826), .CO(n3827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i3 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_41/i2  (.I0(\la0_probe6[1] ), .I1(\la0_probe6[0] ), 
            .CI(1'b0), .O(n3828), .CO(n3829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(297)
    defparam \MCsiRxController/add_41/i2 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_41/i2 .I1_POLARITY = 1'b1;
    EFX_RAM10 \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo  (.WCLK(oTestPort[17]), 
            .RCLK(iSCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd }), 
            .WDATA({\la0_probe9[1] , \la0_probe9[0] , \la0_probe8[7] , 
            \la0_probe8[6] , \la0_probe8[5] , \la0_probe8[4] , \la0_probe8[3] , 
            \la0_probe8[2] , \la0_probe8[1] , \la0_probe8[0] }), .WADDR({\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] }), 
            .RADDR({\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] }), 
            .RDATA({\MCsiRxController/MCsi2Decoder/wFtiRd[9] , \MCsiRxController/MCsi2Decoder/wFtiRd[8] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[7] , \MCsiRxController/MCsi2Decoder/wFtiRd[6] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[5] , \MCsiRxController/MCsi2Decoder/wFtiRd[4] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[3] , \MCsiRxController/MCsi2Decoder/wFtiRd[2] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[1] , \MCsiRxController/MCsi2Decoder/wFtiRd[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=10, WRITE_WIDTH=10, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .READ_WIDTH = 10;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 10;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo  (.WCLK(oTestPort[17]), 
            .RCLK(iSCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd }), 
            .WDATA({3'b000, \la0_probe3[0] , \la0_probe9[7] , \la0_probe9[6] , 
            \la0_probe9[5] , \la0_probe9[4] , \la0_probe9[3] , \la0_probe9[2] }), 
            .WADDR({\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0] }), 
            .RADDR({\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0] }), 
            .RDATA({Open_0, Open_1, Open_2, \MCsiRxController/MCsi2Decoder/wFtiRd[16] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[15] , \MCsiRxController/MCsi2Decoder/wFtiRd[14] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[13] , \MCsiRxController/MCsi2Decoder/wFtiRd[12] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[11] , \MCsiRxController/MCsi2Decoder/wFtiRd[10] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=10, WRITE_WIDTH=10, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .READ_WIDTH = 10;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 10;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo  (.WCLK(iSCLK), 
            .RCLK(iSCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({\MCsiRxController/wHsValid , \MCsiRxController/wHsValid }), 
            .WDATA({\MCsiRxController/wHsPixel[15] , \MCsiRxController/wHsPixel[14] , 
            \MCsiRxController/wHsPixel[13] , \MCsiRxController/wHsPixel[12] , 
            \MCsiRxController/wHsPixel[11] , \MCsiRxController/wHsPixel[10] , 
            \MCsiRxController/wHsPixel[9] , \MCsiRxController/wHsPixel[8] , 
            \MCsiRxController/wHsPixel[7] , \MCsiRxController/wHsPixel[6] , 
            \MCsiRxController/wHsPixel[5] , \MCsiRxController/wHsPixel[4] , 
            \MCsiRxController/wHsPixel[3] , \MCsiRxController/wHsPixel[2] , 
            \MCsiRxController/wHsPixel[1] , \MCsiRxController/wHsPixel[0] }), 
            .WADDR({\MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] }), .RADDR({\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] }), 
            .RDATA({\wVideoPixel[15] , \wVideoPixel[14] , \wVideoPixel[13] , 
            \wVideoPixel[12] , \wVideoPixel[11] , \wVideoPixel[10] , \wVideoPixel[9] , 
            \wVideoPixel[8] , \wVideoPixel[7] , \wVideoPixel[6] , \wVideoPixel[5] , 
            \wVideoPixel[4] , \wVideoPixel[3] , \wVideoPixel[2] , \wVideoPixel[1] , 
            \wVideoPixel[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=16, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="NONE", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .READ_WIDTH = 16;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WRITE_WIDTH = 16;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WE_POLARITY = 2'b11;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RST_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RESET_RAM = "ASYNC";
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RESET_OUTREG = "NONE";
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .OUTPUT_REG = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WRITE_MODE = "READ_FIRST";
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram  (.WCLK(1'b0), 
            .RCLK(iBCLK), .WCLKE(1'b0), .RE(1'b1), .RST(1'b0), .WADDREN(1'b0), 
            .RADDREN(1'b1), .WE({2'b00}), .WADDR({10'b0000000000}), .RADDR({\MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] , 
            \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] , 
            \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] , 
            \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] , 
            \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] , \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0] , 
            \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] }), .RDATA({\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[7] , 
            \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[6] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[5] , 
            \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[4] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[3] , 
            \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[2] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[1] , 
            \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=8, WRITE_WIDTH=8, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="NONE", INIT_0=256'h1F24AD230422DC211D201B1F1C1E001D001CAD1B041A3419E71838160115C0D6, INIT_1=256'hC0962856005508481041772F1B2E7C2D082CAD2B042A00290028352701262425, INIT_2=256'h007F00F980FEE0FDE09A01DFD0E0C0D660BA06AFA4A3A4A2619D309CE09A0398, INIT_3=256'h0000000000000000000000000000000000000000000000000000104101E20094, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .READ_WIDTH = 8;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WRITE_WIDTH = 8;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RESET_OUTREG = "NONE";
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_0 = 256'h1F24AD230422DC211D201B1F1C1E001D001CAD1B041A3419E71838160115C0D6;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1 = 256'hC0962856005508481041772F1B2E7C2D082CAD2B042A00290028352701262425;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_2 = 256'h007F00F980FEE0FDE09A01DFD0E0C0D660BA06AFA4A3A4A2619D309CE09A0398;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000104101E20094;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .OUTPUT_REG = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_SRL8 \MVideoPostProcess/mVideoTimingGen/dff_27/i4_2  (.D(\MVideoPostProcess/mVideoTimingGen/qVrange ), 
            .CLK(iVCLK), .CE(1'b1), .Q(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1 */ ;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_2 .INIT = 8'h0;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_2 .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \MVideoPostProcess/mVideoTimingGen/dff_11/i4_2  (.D(\MVideoPostProcess/mVideoTimingGen/qHrange ), 
            .CLK(iVCLK), .CE(1'b1), .Q(\MVideoPostProcess/mVideoTimingGen/dff_11/i4_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1 */ ;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_2 .INIT = 8'h0;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_2 .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_2 .CE_POLARITY = 1'b1;
    EFX_RAM10 \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[0] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[8]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[1] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[9]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[2] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[10]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[3] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[11]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[4] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[12]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[5] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[13]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[6] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[14]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[7] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[15]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[8] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[0]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[9] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[1]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[10] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[2]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[11] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[3]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[12] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[4]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[13] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[5]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[14] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[6]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[15] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[7]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_LUT4 \edb_top_inst/LUT__3985  (.I0(\edb_top_inst/la0/crc_data_out[17] ), 
            .I1(\edb_top_inst/edb_user_dr[67] ), .I2(\edb_top_inst/la0/crc_data_out[18] ), 
            .I3(\edb_top_inst/edb_user_dr[68] ), .O(\edb_top_inst/n2759 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3985 .LUTMASK = 16'h9009;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[2] , \edb_top_inst/la0/la_biu_inst/fifo_dout[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] }), 
            .WADDR({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i40_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i40_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i40_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i40_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i40_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_2  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_2  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i35_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i35_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i35_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i35_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i35_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i36_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i36_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i36_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i36_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i36_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i37_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i37_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i37_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i37_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i37_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i38_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i38_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i38_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i38_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i38_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i39_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i39_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i39_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i39_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i39_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_2 .CE_POLARITY = 1'b1;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[4] , \edb_top_inst/la0/la_biu_inst/fifo_dout[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[6] , \edb_top_inst/la0/la_biu_inst/fifo_dout[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[8] , \edb_top_inst/la0/la_biu_inst/fifo_dout[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[10] , \edb_top_inst/la0/la_biu_inst/fifo_dout[9] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[12] , \edb_top_inst/la0/la_biu_inst/fifo_dout[11] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[14] , \edb_top_inst/la0/la_biu_inst/fifo_dout[13] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[16] , \edb_top_inst/la0/la_biu_inst/fifo_dout[15] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[18] , \edb_top_inst/la0/la_biu_inst/fifo_dout[17] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[20] , \edb_top_inst/la0/la_biu_inst/fifo_dout[19] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[22] , \edb_top_inst/la0/la_biu_inst/fifo_dout[21] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[24] , \edb_top_inst/la0/la_biu_inst/fifo_dout[23] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[26] , \edb_top_inst/la0/la_biu_inst/fifo_dout[25] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[28] , \edb_top_inst/la0/la_biu_inst/fifo_dout[27] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[30] , \edb_top_inst/la0/la_biu_inst/fifo_dout[29] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[32] , \edb_top_inst/la0/la_biu_inst/fifo_dout[31] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[34] , \edb_top_inst/la0/la_biu_inst/fifo_dout[33] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[36] , \edb_top_inst/la0/la_biu_inst/fifo_dout[35] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[38] , \edb_top_inst/la0/la_biu_inst/fifo_dout[37] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[40] , \edb_top_inst/la0/la_biu_inst/fifo_dout[39] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[42] , \edb_top_inst/la0/la_biu_inst/fifo_dout[41] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_LUT4 \edb_top_inst/LUT__3986  (.I0(\edb_top_inst/la0/crc_data_out[19] ), 
            .I1(\edb_top_inst/edb_user_dr[69] ), .I2(\edb_top_inst/la0/crc_data_out[20] ), 
            .I3(\edb_top_inst/edb_user_dr[70] ), .O(\edb_top_inst/n2760 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3986 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3987  (.I0(\edb_top_inst/la0/crc_data_out[16] ), 
            .I1(\edb_top_inst/edb_user_dr[66] ), .I2(\edb_top_inst/la0/crc_data_out[23] ), 
            .I3(\edb_top_inst/edb_user_dr[73] ), .O(\edb_top_inst/n2761 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3987 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3988  (.I0(\edb_top_inst/n2758 ), .I1(\edb_top_inst/n2759 ), 
            .I2(\edb_top_inst/n2760 ), .I3(\edb_top_inst/n2761 ), .O(\edb_top_inst/n2762 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3988 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3989  (.I0(\edb_top_inst/la0/crc_data_out[24] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/la0/crc_data_out[31] ), 
            .I3(\edb_top_inst/edb_user_dr[81] ), .O(\edb_top_inst/n2763 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3989 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3990  (.I0(\edb_top_inst/la0/crc_data_out[25] ), 
            .I1(\edb_top_inst/edb_user_dr[75] ), .I2(\edb_top_inst/la0/crc_data_out[26] ), 
            .I3(\edb_top_inst/edb_user_dr[76] ), .O(\edb_top_inst/n2764 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3990 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3991  (.I0(\edb_top_inst/la0/crc_data_out[29] ), 
            .I1(\edb_top_inst/edb_user_dr[79] ), .I2(\edb_top_inst/la0/crc_data_out[30] ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n2765 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3991 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3992  (.I0(\edb_top_inst/la0/crc_data_out[27] ), 
            .I1(\edb_top_inst/edb_user_dr[77] ), .I2(\edb_top_inst/la0/crc_data_out[28] ), 
            .I3(\edb_top_inst/edb_user_dr[78] ), .O(\edb_top_inst/n2766 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3992 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3993  (.I0(\edb_top_inst/n2763 ), .I1(\edb_top_inst/n2764 ), 
            .I2(\edb_top_inst/n2765 ), .I3(\edb_top_inst/n2766 ), .O(\edb_top_inst/n2767 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3993 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3994  (.I0(\edb_top_inst/la0/crc_data_out[0] ), 
            .I1(\edb_top_inst/edb_user_dr[50] ), .I2(\edb_top_inst/la0/crc_data_out[1] ), 
            .I3(\edb_top_inst/edb_user_dr[51] ), .O(\edb_top_inst/n2768 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3994 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3995  (.I0(\edb_top_inst/la0/crc_data_out[6] ), 
            .I1(\edb_top_inst/edb_user_dr[56] ), .I2(\edb_top_inst/la0/crc_data_out[15] ), 
            .I3(\edb_top_inst/edb_user_dr[65] ), .O(\edb_top_inst/n2769 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3995 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3996  (.I0(\edb_top_inst/la0/crc_data_out[4] ), 
            .I1(\edb_top_inst/edb_user_dr[54] ), .I2(\edb_top_inst/la0/crc_data_out[5] ), 
            .I3(\edb_top_inst/edb_user_dr[55] ), .O(\edb_top_inst/n2770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3996 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3997  (.I0(\edb_top_inst/la0/crc_data_out[2] ), 
            .I1(\edb_top_inst/edb_user_dr[52] ), .I2(\edb_top_inst/la0/crc_data_out[3] ), 
            .I3(\edb_top_inst/edb_user_dr[53] ), .O(\edb_top_inst/n2771 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3997 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3998  (.I0(\edb_top_inst/n2768 ), .I1(\edb_top_inst/n2769 ), 
            .I2(\edb_top_inst/n2770 ), .I3(\edb_top_inst/n2771 ), .O(\edb_top_inst/n2772 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3998 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3999  (.I0(\edb_top_inst/la0/crc_data_out[8] ), 
            .I1(\edb_top_inst/edb_user_dr[58] ), .I2(\edb_top_inst/la0/crc_data_out[9] ), 
            .I3(\edb_top_inst/edb_user_dr[59] ), .O(\edb_top_inst/n2773 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3999 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4000  (.I0(\edb_top_inst/la0/crc_data_out[10] ), 
            .I1(\edb_top_inst/edb_user_dr[60] ), .I2(\edb_top_inst/la0/crc_data_out[11] ), 
            .I3(\edb_top_inst/edb_user_dr[61] ), .O(\edb_top_inst/n2774 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4000 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4001  (.I0(\edb_top_inst/la0/crc_data_out[12] ), 
            .I1(\edb_top_inst/edb_user_dr[62] ), .I2(\edb_top_inst/la0/crc_data_out[13] ), 
            .I3(\edb_top_inst/edb_user_dr[63] ), .O(\edb_top_inst/n2775 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4001 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4002  (.I0(\edb_top_inst/la0/crc_data_out[7] ), 
            .I1(\edb_top_inst/edb_user_dr[57] ), .I2(\edb_top_inst/la0/crc_data_out[14] ), 
            .I3(\edb_top_inst/edb_user_dr[64] ), .O(\edb_top_inst/n2776 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4002 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4003  (.I0(\edb_top_inst/n2773 ), .I1(\edb_top_inst/n2774 ), 
            .I2(\edb_top_inst/n2775 ), .I3(\edb_top_inst/n2776 ), .O(\edb_top_inst/n2777 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4003 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4004  (.I0(\edb_top_inst/n2762 ), .I1(\edb_top_inst/n2767 ), 
            .I2(\edb_top_inst/n2772 ), .I3(\edb_top_inst/n2777 ), .O(\edb_top_inst/n2778 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4004 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4005  (.I0(\edb_top_inst/la0/bit_count[2] ), 
            .I1(\edb_top_inst/la0/bit_count[3] ), .I2(\edb_top_inst/la0/bit_count[4] ), 
            .I3(\edb_top_inst/la0/bit_count[5] ), .O(\edb_top_inst/n2779 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4005 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4006  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/la0/bit_count[1] ), .I2(\edb_top_inst/n2779 ), 
            .O(\edb_top_inst/n2780 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4006 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4007  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/n2780 ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n2781 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4007 .LUTMASK = 16'h00bf;
    EFX_LUT4 \edb_top_inst/LUT__4008  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n2782 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4008 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4009  (.I0(\edb_top_inst/n2781 ), .I1(\edb_top_inst/n2782 ), 
            .O(\edb_top_inst/n2783 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4009 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4010  (.I0(\edb_top_inst/la0/biu_ready ), 
            .I1(\edb_top_inst/n2778 ), .I2(\edb_top_inst/n2783 ), .O(\edb_top_inst/n2784 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4010 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4011  (.I0(\edb_top_inst/la0/data_out_shift_reg[0] ), 
            .I1(\edb_top_inst/la0/crc_data_out[0] ), .I2(\edb_top_inst/n2783 ), 
            .O(\edb_top_inst/n2785 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4011 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4012  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/n2780 ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n2786 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4012 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__4013  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/n2786 ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .I3(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n2787 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4013 .LUTMASK = 16'h0a0c;
    EFX_LUT4 \edb_top_inst/LUT__4014  (.I0(\edb_top_inst/debug_hub_inst/module_id_reg[1] ), 
            .I1(\edb_top_inst/debug_hub_inst/module_id_reg[2] ), .I2(\edb_top_inst/debug_hub_inst/module_id_reg[3] ), 
            .I3(\edb_top_inst/debug_hub_inst/module_id_reg[0] ), .O(\edb_top_inst/n2788 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4014 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4015  (.I0(\edb_top_inst/n2785 ), .I1(\edb_top_inst/n2784 ), 
            .I2(\edb_top_inst/n2787 ), .I3(\edb_top_inst/n2788 ), .O(jtag_inst2_TDO)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4015 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4016  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[40] ), .O(\edb_top_inst/la0/n1340 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4016 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4017  (.I0(\edb_top_inst/edb_user_dr[81] ), 
            .I1(jtag_inst2_UPDATE), .I2(\edb_top_inst/n2788 ), .O(\edb_top_inst/n2789 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4017 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4018  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n2790 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4018 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4019  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[3] ), .I2(\edb_top_inst/n2790 ), 
            .O(\edb_top_inst/n2791 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4019 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4020  (.I0(\edb_top_inst/edb_user_dr[67] ), 
            .I1(\edb_top_inst/edb_user_dr[68] ), .I2(\edb_top_inst/edb_user_dr[69] ), 
            .I3(\edb_top_inst/edb_user_dr[79] ), .O(\edb_top_inst/n2792 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4020 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4021  (.I0(\edb_top_inst/edb_user_dr[78] ), 
            .I1(\edb_top_inst/edb_user_dr[77] ), .I2(\edb_top_inst/edb_user_dr[80] ), 
            .O(\edb_top_inst/n2793 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4021 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4022  (.I0(\edb_top_inst/n2789 ), .I1(\edb_top_inst/n2791 ), 
            .I2(\edb_top_inst/n2792 ), .I3(\edb_top_inst/n2793 ), .O(\edb_top_inst/n2794 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4022 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4023  (.I0(\edb_top_inst/edb_user_dr[66] ), 
            .I1(\edb_top_inst/n2794 ), .O(\edb_top_inst/n2795 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4023 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4024  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/n2795 ), 
            .O(\edb_top_inst/n2796 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4024 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4025  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .O(\edb_top_inst/n2797 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4025 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4026  (.I0(\edb_top_inst/edb_user_dr[75] ), 
            .I1(\edb_top_inst/edb_user_dr[76] ), .O(\edb_top_inst/n2798 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4026 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4027  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/n2797 ), 
            .I3(\edb_top_inst/n2798 ), .O(\edb_top_inst/n2799 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4027 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4028  (.I0(\edb_top_inst/n2796 ), .I1(\edb_top_inst/n2799 ), 
            .O(\edb_top_inst/la0/n1312 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4028 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4029  (.I0(\edb_top_inst/la0/n1312 ), .I1(\edb_top_inst/la0/la_soft_reset_in ), 
            .O(\edb_top_inst/ceg_net5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4029 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4030  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[41] ), .O(\edb_top_inst/la0/n1341 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4030 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4031  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[42] ), .O(\edb_top_inst/la0/n1342 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4031 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4032  (.I0(\edb_top_inst/edb_user_dr[65] ), 
            .I1(\edb_top_inst/edb_user_dr[64] ), .I2(\edb_top_inst/n2795 ), 
            .O(\edb_top_inst/n2800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4032 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4033  (.I0(\edb_top_inst/n2800 ), .I1(\edb_top_inst/n2799 ), 
            .O(\edb_top_inst/la0/n1396 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4033 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4034  (.I0(\edb_top_inst/n2795 ), .I1(\edb_top_inst/n2799 ), 
            .I2(\edb_top_inst/edb_user_dr[64] ), .I3(\edb_top_inst/edb_user_dr[65] ), 
            .O(\edb_top_inst/la0/n1913 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4034 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4035  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/edb_user_dr[63] ), 
            .I3(\edb_top_inst/edb_user_dr[66] ), .O(\edb_top_inst/n2801 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4035 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4036  (.I0(\edb_top_inst/n2794 ), .I1(\edb_top_inst/n2799 ), 
            .I2(\edb_top_inst/n2801 ), .O(\edb_top_inst/la0/n1965 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4036 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4037  (.I0(\edb_top_inst/la0/address_counter[4] ), 
            .I1(\edb_top_inst/la0/address_counter[5] ), .I2(\edb_top_inst/la0/address_counter[6] ), 
            .I3(\edb_top_inst/la0/address_counter[7] ), .O(\edb_top_inst/n2802 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4037 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4038  (.I0(\edb_top_inst/la0/address_counter[0] ), 
            .I1(\edb_top_inst/la0/address_counter[1] ), .I2(\edb_top_inst/la0/address_counter[2] ), 
            .I3(\edb_top_inst/n2802 ), .O(\edb_top_inst/n2803 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4038 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4039  (.I0(\edb_top_inst/la0/address_counter[8] ), 
            .I1(\edb_top_inst/la0/address_counter[9] ), .I2(\edb_top_inst/la0/address_counter[10] ), 
            .I3(\edb_top_inst/la0/address_counter[11] ), .O(\edb_top_inst/n2804 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4039 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4040  (.I0(\edb_top_inst/la0/address_counter[3] ), 
            .I1(\edb_top_inst/la0/address_counter[12] ), .I2(\edb_top_inst/la0/address_counter[13] ), 
            .I3(\edb_top_inst/la0/address_counter[14] ), .O(\edb_top_inst/n2805 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4040 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4041  (.I0(\edb_top_inst/n2803 ), .I1(\edb_top_inst/n2804 ), 
            .I2(\edb_top_inst/n2805 ), .O(\edb_top_inst/n2806 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4041 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4042  (.I0(\edb_top_inst/n2806 ), .I1(\edb_top_inst/n67 ), 
            .I2(\edb_top_inst/edb_user_dr[45] ), .I3(\edb_top_inst/n2791 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4042 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4043  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/la0/module_state[2] ), 
            .I2(\edb_top_inst/la0/module_state[3] ), .I3(\edb_top_inst/la0/biu_ready ), 
            .O(\edb_top_inst/n2807 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4043 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4044  (.I0(\edb_top_inst/n2807 ), .I1(\edb_top_inst/la0/module_state[0] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n2808 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4044 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4045  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[2] ), 
            .I3(\edb_top_inst/la0/word_count[3] ), .O(\edb_top_inst/n2809 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4045 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4046  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/la0/word_count[6] ), 
            .I3(\edb_top_inst/n2809 ), .O(\edb_top_inst/n2810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4046 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4047  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n2811 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4047 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4048  (.I0(\edb_top_inst/la0/word_count[1] ), 
            .I1(\edb_top_inst/la0/word_count[2] ), .I2(\edb_top_inst/la0/word_count[7] ), 
            .I3(\edb_top_inst/la0/word_count[8] ), .O(\edb_top_inst/n2812 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4048 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4049  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/la0/word_count[14] ), 
            .I3(\edb_top_inst/n2812 ), .O(\edb_top_inst/n2813 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4049 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4050  (.I0(\edb_top_inst/la0/word_count[9] ), 
            .I1(\edb_top_inst/la0/word_count[10] ), .I2(\edb_top_inst/la0/word_count[11] ), 
            .I3(\edb_top_inst/la0/word_count[12] ), .O(\edb_top_inst/n2814 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4050 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4051  (.I0(\edb_top_inst/la0/word_count[3] ), 
            .I1(\edb_top_inst/la0/word_count[6] ), .I2(\edb_top_inst/la0/word_count[13] ), 
            .I3(\edb_top_inst/la0/word_count[15] ), .O(\edb_top_inst/n2815 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4051 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4052  (.I0(\edb_top_inst/n2813 ), .I1(\edb_top_inst/n2814 ), 
            .I2(\edb_top_inst/n2815 ), .O(\edb_top_inst/n2816 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4052 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4053  (.I0(\edb_top_inst/n2810 ), .I1(\edb_top_inst/n2808 ), 
            .I2(\edb_top_inst/n2816 ), .I3(\edb_top_inst/n2811 ), .O(\edb_top_inst/n2817 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5f0c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4053 .LUTMASK = 16'h5f0c;
    EFX_LUT4 \edb_top_inst/LUT__4054  (.I0(\edb_top_inst/n2790 ), .I1(\edb_top_inst/n2817 ), 
            .I2(\edb_top_inst/la0/module_state[2] ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n2818 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4054 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__4055  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/n2819 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4055 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__4056  (.I0(\edb_top_inst/n2819 ), .I1(\edb_top_inst/la0/bit_count[0] ), 
            .I2(\edb_top_inst/la0/bit_count[1] ), .I3(\edb_top_inst/la0/bit_count[2] ), 
            .O(\edb_top_inst/n2820 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbffd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4056 .LUTMASK = 16'hbffd;
    EFX_LUT4 \edb_top_inst/LUT__4057  (.I0(\edb_top_inst/la0/opcode[3] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[0] ), .O(\edb_top_inst/n2736 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4057 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4058  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/n2733 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4058 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4059  (.I0(\edb_top_inst/n2736 ), .I1(\edb_top_inst/n2733 ), 
            .I2(\edb_top_inst/la0/bit_count[5] ), .I3(\edb_top_inst/la0/bit_count[4] ), 
            .O(\edb_top_inst/n2821 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3dfe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4059 .LUTMASK = 16'h3dfe;
    EFX_LUT4 \edb_top_inst/LUT__4060  (.I0(\edb_top_inst/la0/opcode[1] ), 
            .I1(\edb_top_inst/la0/opcode[3] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[0] ), .O(\edb_top_inst/n1249 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4060 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4061  (.I0(\edb_top_inst/n2819 ), .I1(\edb_top_inst/n1249 ), 
            .O(\edb_top_inst/n2822 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4061 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4062  (.I0(\edb_top_inst/n2820 ), .I1(\edb_top_inst/n2821 ), 
            .I2(\edb_top_inst/n2822 ), .I3(\edb_top_inst/la0/bit_count[3] ), 
            .O(\edb_top_inst/n2823 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4062 .LUTMASK = 16'h1001;
    EFX_LUT4 \edb_top_inst/LUT__4063  (.I0(\edb_top_inst/n2816 ), .I1(\edb_top_inst/la0/module_state[0] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/n2823 ), 
            .O(\edb_top_inst/n2824 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4063 .LUTMASK = 16'hc100;
    EFX_LUT4 \edb_top_inst/LUT__4064  (.I0(\edb_top_inst/n2824 ), .I1(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n2825 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4064 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4065  (.I0(\edb_top_inst/edb_user_dr[77] ), 
            .I1(\edb_top_inst/edb_user_dr[78] ), .I2(\edb_top_inst/edb_user_dr[79] ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n2826 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4065 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__4066  (.I0(\edb_top_inst/n2826 ), .I1(\edb_top_inst/la0/module_state[2] ), 
            .I2(\edb_top_inst/n2789 ), .I3(\edb_top_inst/n2790 ), .O(\edb_top_inst/n2827 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4066 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4067  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/n2827 ), .O(\edb_top_inst/la0/op_reg_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4067 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4068  (.I0(\edb_top_inst/n2825 ), .I1(\edb_top_inst/n2818 ), 
            .I2(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/addr_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4068 .LUTMASK = 16'hf4f4;
    EFX_LUT4 \edb_top_inst/LUT__4069  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/la0/module_state[2] ), .O(\edb_top_inst/n2828 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4069 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4070  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/n2823 ), 
            .I3(\edb_top_inst/n2828 ), .O(\edb_top_inst/n2829 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4070 .LUTMASK = 16'h9000;
    EFX_LUT4 \edb_top_inst/LUT__4071  (.I0(\edb_top_inst/n2782 ), .I1(\edb_top_inst/n2790 ), 
            .O(\edb_top_inst/n2830 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4071 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4072  (.I0(\edb_top_inst/n2829 ), .I1(\edb_top_inst/n2827 ), 
            .I2(\edb_top_inst/n2808 ), .I3(\edb_top_inst/n2830 ), .O(\edb_top_inst/n2831 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4072 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4073  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/n2831 ), .O(\edb_top_inst/la0/n2189 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4073 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4074  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n2832 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4074 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4075  (.I0(\edb_top_inst/edb_user_dr[81] ), 
            .I1(\edb_top_inst/n2832 ), .I2(\edb_top_inst/n2788 ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n2833 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4075 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__4076  (.I0(\edb_top_inst/n2833 ), .I1(\edb_top_inst/la0/module_state[0] ), 
            .I2(\edb_top_inst/n2828 ), .O(\edb_top_inst/n2834 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4076 .LUTMASK = 16'h9090;
    EFX_LUT4 \edb_top_inst/LUT__4077  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/n2782 ), .I2(\edb_top_inst/n2834 ), .I3(\edb_top_inst/n2831 ), 
            .O(\edb_top_inst/ceg_net26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4077 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__4078  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/edb_user_dr[29] ), .I2(\edb_top_inst/n2791 ), 
            .O(\edb_top_inst/la0/data_to_word_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4078 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4079  (.I0(\edb_top_inst/n2816 ), .I1(\edb_top_inst/n2810 ), 
            .O(\edb_top_inst/n2835 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4079 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4080  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n2836 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4080 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4081  (.I0(\edb_top_inst/n2823 ), .I1(\edb_top_inst/n2835 ), 
            .I2(\edb_top_inst/n2836 ), .I3(\edb_top_inst/n2833 ), .O(\edb_top_inst/n2837 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4081 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__4082  (.I0(\edb_top_inst/n2816 ), .I1(\edb_top_inst/n2810 ), 
            .I2(\edb_top_inst/n2832 ), .O(\edb_top_inst/n2838 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4082 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4083  (.I0(\edb_top_inst/n2788 ), .I1(jtag_inst2_CAPTURE), 
            .O(\edb_top_inst/n2839 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4083 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4084  (.I0(\edb_top_inst/n2810 ), .I1(\edb_top_inst/n2816 ), 
            .I2(\edb_top_inst/n2839 ), .I3(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n2840 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4084 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__4085  (.I0(\edb_top_inst/n2823 ), .I1(\edb_top_inst/n2838 ), 
            .I2(\edb_top_inst/n2840 ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n2841 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4085 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4086  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/la0/biu_ready ), 
            .I2(\edb_top_inst/n2839 ), .I3(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n2842 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4086 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4087  (.I0(\edb_top_inst/n2842 ), .I1(\edb_top_inst/la0/module_state[2] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/n2827 ), 
            .O(\edb_top_inst/n2843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4087 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__4088  (.I0(\edb_top_inst/n2841 ), .I1(\edb_top_inst/n2837 ), 
            .I2(\edb_top_inst/la0/module_state[2] ), .I3(\edb_top_inst/n2843 ), 
            .O(\edb_top_inst/n2844 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4088 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__4089  (.I0(\edb_top_inst/n2844 ), .I1(\edb_top_inst/la0/module_state[0] ), 
            .I2(\edb_top_inst/n2828 ), .I3(\edb_top_inst/n2831 ), .O(\edb_top_inst/la0/word_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h10ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4089 .LUTMASK = 16'h10ff;
    EFX_LUT4 \edb_top_inst/LUT__4090  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/n2845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hec07, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4090 .LUTMASK = 16'hec07;
    EFX_LUT4 \edb_top_inst/LUT__4091  (.I0(\edb_top_inst/la0/internal_register_select[10] ), 
            .I1(\edb_top_inst/la0/internal_register_select[11] ), .I2(\edb_top_inst/la0/internal_register_select[12] ), 
            .O(\edb_top_inst/n2846 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4091 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4092  (.I0(\edb_top_inst/la0/internal_register_select[1] ), 
            .I1(\edb_top_inst/la0/internal_register_select[2] ), .I2(\edb_top_inst/la0/internal_register_select[4] ), 
            .I3(\edb_top_inst/la0/internal_register_select[5] ), .O(\edb_top_inst/n2847 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4092 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4093  (.I0(\edb_top_inst/la0/internal_register_select[6] ), 
            .I1(\edb_top_inst/la0/internal_register_select[7] ), .I2(\edb_top_inst/la0/internal_register_select[8] ), 
            .I3(\edb_top_inst/la0/internal_register_select[9] ), .O(\edb_top_inst/n2848 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4093 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4094  (.I0(\edb_top_inst/n2846 ), .I1(\edb_top_inst/n2847 ), 
            .I2(\edb_top_inst/n2848 ), .O(\edb_top_inst/n2849 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4094 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4095  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/n2849 ), .O(\edb_top_inst/n2850 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4095 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4096  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4096 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4097  (.I0(\edb_top_inst/n2849 ), .I1(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n2852 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4097 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4098  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/n2852 ), .O(\edb_top_inst/n2853 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4098 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4099  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[0] ), 
            .I2(\edb_top_inst/n2845 ), .I3(\edb_top_inst/n2851 ), .O(\edb_top_inst/n2854 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4099 .LUTMASK = 16'h7077;
    EFX_LUT4 \edb_top_inst/LUT__4100  (.I0(\edb_top_inst/n2828 ), .I1(\edb_top_inst/n2823 ), 
            .I2(\edb_top_inst/n2790 ), .I3(\edb_top_inst/n2808 ), .O(\edb_top_inst/n2855 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4100 .LUTMASK = 16'h007f;
    EFX_LUT4 \edb_top_inst/LUT__4101  (.I0(\edb_top_inst/la0/data_from_biu[0] ), 
            .I1(\edb_top_inst/n2854 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2856 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4101 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4102  (.I0(\edb_top_inst/n2839 ), .I1(\edb_top_inst/n2791 ), 
            .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2857 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4102 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__4103  (.I0(\edb_top_inst/la0/data_out_shift_reg[1] ), 
            .I1(\edb_top_inst/n2856 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4103 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4104  (.I0(jtag_inst2_CAPTURE), .I1(jtag_inst2_SHIFT), 
            .I2(\edb_top_inst/n2788 ), .I3(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n2858 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4104 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__4105  (.I0(\edb_top_inst/n2858 ), .I1(\edb_top_inst/la0/module_state[3] ), 
            .I2(\edb_top_inst/n2790 ), .I3(\edb_top_inst/n2808 ), .O(\edb_top_inst/ceg_net14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4105 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__4106  (.I0(\edb_top_inst/n2780 ), .I1(\edb_top_inst/n2835 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n2859 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4106 .LUTMASK = 16'h050c;
    EFX_LUT4 \edb_top_inst/LUT__4107  (.I0(\edb_top_inst/n2859 ), .I1(jtag_inst2_UPDATE), 
            .I2(\edb_top_inst/la0/module_state[2] ), .O(\edb_top_inst/n2860 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4107 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4108  (.I0(\edb_top_inst/n2860 ), .I1(\edb_top_inst/n2844 ), 
            .I2(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/la0/module_next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4108 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__4109  (.I0(\edb_top_inst/edb_user_dr[74] ), 
            .I1(\edb_top_inst/edb_user_dr[73] ), .I2(\edb_top_inst/n2798 ), 
            .O(\edb_top_inst/n2861 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4109 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4110  (.I0(\edb_top_inst/n2861 ), .I1(\edb_top_inst/n2797 ), 
            .O(\edb_top_inst/n2862 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4110 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4111  (.I0(\edb_top_inst/n2800 ), .I1(\edb_top_inst/n2862 ), 
            .O(\edb_top_inst/la0/n5294 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4111 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4112  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/n2795 ), .I2(\edb_top_inst/edb_user_dr[65] ), 
            .O(\edb_top_inst/n2863 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4112 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4113  (.I0(\edb_top_inst/n2863 ), .I1(\edb_top_inst/n2862 ), 
            .O(\edb_top_inst/la0/n5492 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4113 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4114  (.I0(\edb_top_inst/n2796 ), .I1(\edb_top_inst/n2861 ), 
            .O(\edb_top_inst/n2864 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4114 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4115  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .O(\edb_top_inst/n2865 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4115 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4116  (.I0(\edb_top_inst/n2864 ), .I1(\edb_top_inst/n2865 ), 
            .O(\edb_top_inst/la0/n6947 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4116 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4117  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/n2861 ), .I2(\edb_top_inst/edb_user_dr[71] ), 
            .I3(\edb_top_inst/edb_user_dr[72] ), .O(\edb_top_inst/n2866 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4117 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4118  (.I0(\edb_top_inst/n2800 ), .I1(\edb_top_inst/n2866 ), 
            .O(\edb_top_inst/la0/n7907 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4118 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4119  (.I0(\edb_top_inst/n2863 ), .I1(\edb_top_inst/n2866 ), 
            .O(\edb_top_inst/la0/n8105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4119 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4120  (.I0(\edb_top_inst/n2798 ), .I1(\edb_top_inst/edb_user_dr[74] ), 
            .O(\edb_top_inst/n2867 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4120 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4121  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/n2867 ), .O(\edb_top_inst/n2868 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4121 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4122  (.I0(\edb_top_inst/n2796 ), .I1(\edb_top_inst/n2868 ), 
            .O(\edb_top_inst/n2869 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4122 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4123  (.I0(\edb_top_inst/n2869 ), .I1(\edb_top_inst/n2797 ), 
            .O(\edb_top_inst/la0/n8741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4123 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4124  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[72] ), .I2(\edb_top_inst/edb_user_dr[71] ), 
            .O(\edb_top_inst/n2870 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4124 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4125  (.I0(\edb_top_inst/n2800 ), .I1(\edb_top_inst/n2868 ), 
            .I2(\edb_top_inst/n2870 ), .O(\edb_top_inst/la0/n9645 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4125 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4126  (.I0(\edb_top_inst/n2863 ), .I1(\edb_top_inst/n2868 ), 
            .I2(\edb_top_inst/n2870 ), .O(\edb_top_inst/la0/n9843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4126 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4127  (.I0(\edb_top_inst/n2869 ), .I1(\edb_top_inst/n2865 ), 
            .O(\edb_top_inst/la0/n10527 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4127 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4128  (.I0(\edb_top_inst/n2800 ), .I1(\edb_top_inst/n2868 ), 
            .I2(\edb_top_inst/n2865 ), .O(\edb_top_inst/la0/n10542 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4128 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4129  (.I0(\edb_top_inst/n2863 ), .I1(\edb_top_inst/n2868 ), 
            .I2(\edb_top_inst/n2865 ), .O(\edb_top_inst/la0/n10740 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4129 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4130  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/n2869 ), .I2(\edb_top_inst/edb_user_dr[71] ), 
            .I3(\edb_top_inst/edb_user_dr[72] ), .O(\edb_top_inst/la0/n11368 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4130 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4131  (.I0(\edb_top_inst/n2796 ), .I1(\edb_top_inst/n2867 ), 
            .I2(\edb_top_inst/n2797 ), .I3(\edb_top_inst/edb_user_dr[73] ), 
            .O(\edb_top_inst/la0/n12201 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4131 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4132  (.I0(\edb_top_inst/n2789 ), .I1(\edb_top_inst/n2791 ), 
            .I2(\edb_top_inst/n2793 ), .O(\edb_top_inst/la0/regsel_ld_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4132 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4133  (.I0(\edb_top_inst/n2806 ), .I1(\edb_top_inst/n1112 ), 
            .I2(\edb_top_inst/edb_user_dr[46] ), .I3(\edb_top_inst/n2791 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4133 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4134  (.I0(\edb_top_inst/n2806 ), .I1(\edb_top_inst/n1110 ), 
            .I2(\edb_top_inst/edb_user_dr[47] ), .I3(\edb_top_inst/n2791 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4134 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4135  (.I0(\edb_top_inst/n2806 ), .I1(\edb_top_inst/n1108 ), 
            .I2(\edb_top_inst/edb_user_dr[48] ), .I3(\edb_top_inst/n2791 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4135 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4136  (.I0(\edb_top_inst/n1106 ), .I1(\edb_top_inst/edb_user_dr[49] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4136 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4137  (.I0(\edb_top_inst/n1104 ), .I1(\edb_top_inst/edb_user_dr[50] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4137 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4138  (.I0(\edb_top_inst/n1102 ), .I1(\edb_top_inst/edb_user_dr[51] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4138 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4139  (.I0(\edb_top_inst/n1100 ), .I1(\edb_top_inst/edb_user_dr[52] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4139 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4140  (.I0(\edb_top_inst/n1098 ), .I1(\edb_top_inst/edb_user_dr[53] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4140 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4141  (.I0(\edb_top_inst/n1096 ), .I1(\edb_top_inst/edb_user_dr[54] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4141 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4142  (.I0(\edb_top_inst/n1094 ), .I1(\edb_top_inst/edb_user_dr[55] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4142 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4143  (.I0(\edb_top_inst/n1092 ), .I1(\edb_top_inst/edb_user_dr[56] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4143 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4144  (.I0(\edb_top_inst/n1090 ), .I1(\edb_top_inst/edb_user_dr[57] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4144 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4145  (.I0(\edb_top_inst/n1088 ), .I1(\edb_top_inst/edb_user_dr[58] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4145 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4146  (.I0(\edb_top_inst/n1086 ), .I1(\edb_top_inst/edb_user_dr[59] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4146 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4147  (.I0(\edb_top_inst/n1084 ), .I1(\edb_top_inst/la0/address_counter[15] ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2871 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4147 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4148  (.I0(\edb_top_inst/edb_user_dr[60] ), 
            .I1(\edb_top_inst/n2871 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4148 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4149  (.I0(\edb_top_inst/n1082 ), .I1(\edb_top_inst/n1146 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2872 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4149 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4150  (.I0(\edb_top_inst/edb_user_dr[61] ), 
            .I1(\edb_top_inst/n2872 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4150 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4151  (.I0(\edb_top_inst/n1080 ), .I1(\edb_top_inst/n1144 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2873 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4151 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4152  (.I0(\edb_top_inst/edb_user_dr[62] ), 
            .I1(\edb_top_inst/n2873 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4152 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4153  (.I0(\edb_top_inst/n1078 ), .I1(\edb_top_inst/n1142 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2874 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4153 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4154  (.I0(\edb_top_inst/edb_user_dr[63] ), 
            .I1(\edb_top_inst/n2874 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4154 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4155  (.I0(\edb_top_inst/n1076 ), .I1(\edb_top_inst/n1137 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2875 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4155 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4156  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/n2875 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4156 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4157  (.I0(\edb_top_inst/n1074 ), .I1(\edb_top_inst/n1135 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2876 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4157 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4158  (.I0(\edb_top_inst/edb_user_dr[65] ), 
            .I1(\edb_top_inst/n2876 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4158 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4159  (.I0(\edb_top_inst/n1072 ), .I1(\edb_top_inst/n1133 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2877 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4159 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4160  (.I0(\edb_top_inst/edb_user_dr[66] ), 
            .I1(\edb_top_inst/n2877 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4160 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4161  (.I0(\edb_top_inst/n1070 ), .I1(\edb_top_inst/n1131 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2878 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4161 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4162  (.I0(\edb_top_inst/edb_user_dr[67] ), 
            .I1(\edb_top_inst/n2878 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4162 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4163  (.I0(\edb_top_inst/n1068 ), .I1(\edb_top_inst/n1129 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2879 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4163 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4164  (.I0(\edb_top_inst/edb_user_dr[68] ), 
            .I1(\edb_top_inst/n2879 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4164 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4165  (.I0(\edb_top_inst/n1066 ), .I1(\edb_top_inst/n1127 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2880 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4165 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4166  (.I0(\edb_top_inst/edb_user_dr[69] ), 
            .I1(\edb_top_inst/n2880 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4166 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4167  (.I0(\edb_top_inst/n1064 ), .I1(\edb_top_inst/n1125 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2881 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4167 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4168  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/n2881 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4168 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4169  (.I0(\edb_top_inst/n1062 ), .I1(\edb_top_inst/n1123 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2882 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4169 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4170  (.I0(\edb_top_inst/edb_user_dr[71] ), 
            .I1(\edb_top_inst/n2882 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4170 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4181  (.I0(\edb_top_inst/n2831 ), .I1(\edb_top_inst/n69 ), 
            .O(\edb_top_inst/la0/n2188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4181 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4182  (.I0(\edb_top_inst/n2831 ), .I1(\edb_top_inst/n1051 ), 
            .O(\edb_top_inst/la0/n2187 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4182 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4183  (.I0(\edb_top_inst/n2831 ), .I1(\edb_top_inst/n1049 ), 
            .O(\edb_top_inst/la0/n2186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4183 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4184  (.I0(\edb_top_inst/n2831 ), .I1(\edb_top_inst/n1047 ), 
            .O(\edb_top_inst/la0/n2185 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4184 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4185  (.I0(\edb_top_inst/n2831 ), .I1(\edb_top_inst/n1046 ), 
            .O(\edb_top_inst/la0/n2184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4185 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4186  (.I0(\edb_top_inst/edb_user_dr[30] ), 
            .I1(\edb_top_inst/la0/word_count[0] ), .I2(\edb_top_inst/la0/word_count[1] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haac3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4186 .LUTMASK = 16'haac3;
    EFX_LUT4 \edb_top_inst/LUT__4187  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[2] ), 
            .O(\edb_top_inst/n2888 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he1e1, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4187 .LUTMASK = 16'he1e1;
    EFX_LUT4 \edb_top_inst/LUT__4188  (.I0(\edb_top_inst/n2888 ), .I1(\edb_top_inst/edb_user_dr[31] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4188 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4189  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[2] ), 
            .I3(\edb_top_inst/la0/word_count[3] ), .O(\edb_top_inst/n2889 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe01, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4189 .LUTMASK = 16'hfe01;
    EFX_LUT4 \edb_top_inst/LUT__4190  (.I0(\edb_top_inst/n2889 ), .I1(\edb_top_inst/edb_user_dr[32] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4190 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4191  (.I0(\edb_top_inst/edb_user_dr[33] ), 
            .I1(\edb_top_inst/n2809 ), .I2(\edb_top_inst/la0/word_count[4] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4191 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4192  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/n2809 ), .I2(\edb_top_inst/la0/word_count[5] ), 
            .O(\edb_top_inst/n2890 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4192 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__4193  (.I0(\edb_top_inst/n2890 ), .I1(\edb_top_inst/edb_user_dr[34] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4193 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4194  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/n2809 ), 
            .I3(\edb_top_inst/la0/word_count[6] ), .O(\edb_top_inst/n2891 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4194 .LUTMASK = 16'hef10;
    EFX_LUT4 \edb_top_inst/LUT__4195  (.I0(\edb_top_inst/n2891 ), .I1(\edb_top_inst/edb_user_dr[35] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4195 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4196  (.I0(\edb_top_inst/edb_user_dr[36] ), 
            .I1(\edb_top_inst/n2810 ), .I2(\edb_top_inst/la0/word_count[7] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4196 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4197  (.I0(\edb_top_inst/la0/word_count[7] ), 
            .I1(\edb_top_inst/n2810 ), .I2(\edb_top_inst/la0/word_count[8] ), 
            .O(\edb_top_inst/n2892 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4197 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__4198  (.I0(\edb_top_inst/edb_user_dr[37] ), 
            .I1(\edb_top_inst/n2892 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4198 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4199  (.I0(\edb_top_inst/la0/word_count[7] ), 
            .I1(\edb_top_inst/la0/word_count[8] ), .I2(\edb_top_inst/n2810 ), 
            .O(\edb_top_inst/n2893 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4199 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4200  (.I0(\edb_top_inst/edb_user_dr[38] ), 
            .I1(\edb_top_inst/n2893 ), .I2(\edb_top_inst/la0/word_count[9] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4200 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4201  (.I0(\edb_top_inst/la0/word_count[9] ), 
            .I1(\edb_top_inst/n2893 ), .O(\edb_top_inst/n2894 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4201 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4202  (.I0(\edb_top_inst/edb_user_dr[39] ), 
            .I1(\edb_top_inst/n2894 ), .I2(\edb_top_inst/la0/word_count[10] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4202 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4203  (.I0(\edb_top_inst/la0/word_count[10] ), 
            .I1(\edb_top_inst/n2894 ), .O(\edb_top_inst/n2895 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4203 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4204  (.I0(\edb_top_inst/edb_user_dr[40] ), 
            .I1(\edb_top_inst/n2895 ), .I2(\edb_top_inst/la0/word_count[11] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4204 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4205  (.I0(\edb_top_inst/la0/word_count[11] ), 
            .I1(\edb_top_inst/n2895 ), .O(\edb_top_inst/n2896 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4205 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4206  (.I0(\edb_top_inst/edb_user_dr[41] ), 
            .I1(\edb_top_inst/n2896 ), .I2(\edb_top_inst/la0/word_count[12] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4206 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4207  (.I0(\edb_top_inst/n2893 ), .I1(\edb_top_inst/n2814 ), 
            .O(\edb_top_inst/n2897 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4207 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4208  (.I0(\edb_top_inst/edb_user_dr[42] ), 
            .I1(\edb_top_inst/n2897 ), .I2(\edb_top_inst/la0/word_count[13] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4208 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4209  (.I0(\edb_top_inst/la0/word_count[13] ), 
            .I1(\edb_top_inst/n2897 ), .O(\edb_top_inst/n2898 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4209 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4210  (.I0(\edb_top_inst/edb_user_dr[43] ), 
            .I1(\edb_top_inst/n2898 ), .I2(\edb_top_inst/la0/word_count[14] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4210 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4211  (.I0(\edb_top_inst/la0/word_count[14] ), 
            .I1(\edb_top_inst/n2898 ), .I2(\edb_top_inst/la0/word_count[15] ), 
            .O(\edb_top_inst/n2899 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4211 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__4212  (.I0(\edb_top_inst/edb_user_dr[44] ), 
            .I1(\edb_top_inst/n2899 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4212 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__4213  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2900 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4213 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4214  (.I0(\edb_top_inst/n2851 ), .I1(\edb_top_inst/n2808 ), 
            .I2(\edb_top_inst/n2828 ), .O(\edb_top_inst/n2901 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4214 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4215  (.I0(\edb_top_inst/la0/data_from_biu[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[1] ), .I2(\edb_top_inst/n2900 ), 
            .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2902 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4215 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__4216  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n2903 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4216 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4217  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n2904 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4217 .LUTMASK = 16'hd3d3;
    EFX_LUT4 \edb_top_inst/LUT__4218  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/n2903 ), .I2(\edb_top_inst/n2904 ), .O(\edb_top_inst/n2905 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4218 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4219  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/n2849 ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .O(\edb_top_inst/n2906 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4219 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4220  (.I0(\edb_top_inst/n2851 ), .I1(\edb_top_inst/n2905 ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2907 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4220 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4221  (.I0(\edb_top_inst/n2907 ), .I1(\edb_top_inst/n2902 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[2] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2465 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4221 .LUTMASK = 16'hf0ee;
    EFX_LUT4 \edb_top_inst/LUT__4222  (.I0(\edb_top_inst/la0/data_from_biu[2] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[2] ), .I2(\edb_top_inst/n2900 ), 
            .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2908 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4222 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__4223  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n2909 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4223 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4224  (.I0(\edb_top_inst/n2851 ), .I1(\edb_top_inst/n2909 ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2910 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4224 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4225  (.I0(\edb_top_inst/n2910 ), .I1(\edb_top_inst/n2908 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[3] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2464 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4225 .LUTMASK = 16'hf0ee;
    EFX_LUT4 \edb_top_inst/LUT__4226  (.I0(\edb_top_inst/la0/data_from_biu[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[3] ), .I2(\edb_top_inst/n2900 ), 
            .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2911 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4226 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4227  (.I0(\edb_top_inst/la0/la_sample_cnt[0] ), 
            .I1(\edb_top_inst/la0/internal_register_select[0] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .O(\edb_top_inst/n2912 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3d3d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4227 .LUTMASK = 16'h3d3d;
    EFX_LUT4 \edb_top_inst/LUT__4228  (.I0(\edb_top_inst/n2912 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/n2900 ), .O(\edb_top_inst/n2913 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4228 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4229  (.I0(\edb_top_inst/n2913 ), .I1(\edb_top_inst/n2911 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[4] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2463 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4229 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4230  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[4] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2914 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4230 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4231  (.I0(\edb_top_inst/la0/data_from_biu[4] ), 
            .I1(\edb_top_inst/n2914 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2915 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4231 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4232  (.I0(\edb_top_inst/n2915 ), .I1(\edb_top_inst/la0/data_out_shift_reg[5] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4232 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4233  (.I0(\edb_top_inst/la0/la_sample_cnt[2] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[5] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2916 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4233 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4234  (.I0(\edb_top_inst/la0/data_from_biu[5] ), 
            .I1(\edb_top_inst/n2916 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2917 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4234 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4235  (.I0(\edb_top_inst/n2917 ), .I1(\edb_top_inst/la0/data_out_shift_reg[6] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4235 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4236  (.I0(\edb_top_inst/la0/la_sample_cnt[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[6] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2918 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4236 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4237  (.I0(\edb_top_inst/n2918 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[6] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2919 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4237 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4238  (.I0(\edb_top_inst/n2919 ), .I1(\edb_top_inst/la0/data_out_shift_reg[7] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4238 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4239  (.I0(\edb_top_inst/la0/la_sample_cnt[4] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[7] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2920 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4239 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4240  (.I0(\edb_top_inst/n2920 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[7] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2921 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4240 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4241  (.I0(\edb_top_inst/n2921 ), .I1(\edb_top_inst/la0/data_out_shift_reg[8] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2459 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4241 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4242  (.I0(\edb_top_inst/la0/la_sample_cnt[5] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[8] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2922 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4242 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4243  (.I0(\edb_top_inst/n2922 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[8] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2923 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4243 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4244  (.I0(\edb_top_inst/n2923 ), .I1(\edb_top_inst/la0/data_out_shift_reg[9] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4244 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4245  (.I0(\edb_top_inst/la0/la_sample_cnt[6] ), 
            .I1(\edb_top_inst/n2901 ), .I2(\edb_top_inst/n2852 ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2924 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4245 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4246  (.I0(\edb_top_inst/la0/la_trig_mask[9] ), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/la0/data_from_biu[9] ), 
            .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2925 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4246 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__4247  (.I0(\edb_top_inst/n2924 ), .I1(\edb_top_inst/n2925 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[10] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2457 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4247 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4248  (.I0(\edb_top_inst/la0/la_sample_cnt[7] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[10] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2926 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4248 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4249  (.I0(\edb_top_inst/la0/data_from_biu[10] ), 
            .I1(\edb_top_inst/n2926 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2927 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4249 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4250  (.I0(\edb_top_inst/n2927 ), .I1(\edb_top_inst/la0/data_out_shift_reg[11] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4250 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4251  (.I0(\edb_top_inst/la0/la_sample_cnt[8] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[11] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2928 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4251 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4252  (.I0(\edb_top_inst/n2928 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[11] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2929 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4252 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4253  (.I0(\edb_top_inst/n2929 ), .I1(\edb_top_inst/la0/data_out_shift_reg[12] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2455 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4253 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4254  (.I0(\edb_top_inst/la0/la_sample_cnt[9] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[12] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2930 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4254 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4255  (.I0(\edb_top_inst/n2930 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[12] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2931 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4255 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4256  (.I0(\edb_top_inst/n2931 ), .I1(\edb_top_inst/la0/data_out_shift_reg[13] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4256 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4257  (.I0(\edb_top_inst/la0/la_sample_cnt[10] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[13] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2932 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4257 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4258  (.I0(\edb_top_inst/la0/data_from_biu[13] ), 
            .I1(\edb_top_inst/n2932 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2933 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4258 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4259  (.I0(\edb_top_inst/n2933 ), .I1(\edb_top_inst/la0/data_out_shift_reg[14] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2453 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4259 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4260  (.I0(\edb_top_inst/la0/la_sample_cnt[11] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[14] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2934 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4260 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4261  (.I0(\edb_top_inst/n2934 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[14] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2935 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4261 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4262  (.I0(\edb_top_inst/n2935 ), .I1(\edb_top_inst/la0/data_out_shift_reg[15] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4262 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4263  (.I0(\edb_top_inst/la0/la_sample_cnt[12] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[15] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2936 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4263 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4264  (.I0(\edb_top_inst/n2936 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[15] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2937 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4264 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4265  (.I0(\edb_top_inst/n2937 ), .I1(\edb_top_inst/la0/data_out_shift_reg[16] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4265 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4266  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[16] ), .I2(\edb_top_inst/n2852 ), 
            .O(\edb_top_inst/n2938 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4266 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__4267  (.I0(\edb_top_inst/la0/data_from_biu[16] ), 
            .I1(\edb_top_inst/n2938 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2939 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4267 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4268  (.I0(\edb_top_inst/n2939 ), .I1(\edb_top_inst/la0/data_out_shift_reg[17] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4268 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4269  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[17] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/n2849 ), .O(\edb_top_inst/n2940 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4269 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4270  (.I0(\edb_top_inst/la0/data_from_biu[17] ), 
            .I1(\edb_top_inst/n2940 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2941 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4270 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4271  (.I0(\edb_top_inst/n2941 ), .I1(\edb_top_inst/la0/data_out_shift_reg[18] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2449 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4271 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4272  (.I0(\edb_top_inst/n2850 ), .I1(\edb_top_inst/la0/internal_register_select[0] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[18] ), .O(\edb_top_inst/n2942 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4272 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4273  (.I0(\edb_top_inst/la0/data_from_biu[18] ), 
            .I1(\edb_top_inst/n2942 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2943 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4273 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4274  (.I0(\edb_top_inst/n2943 ), .I1(\edb_top_inst/la0/data_out_shift_reg[19] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4274 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4275  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[19] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/n2849 ), .O(\edb_top_inst/n2944 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4275 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4276  (.I0(\edb_top_inst/la0/data_from_biu[19] ), 
            .I1(\edb_top_inst/n2944 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2945 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4276 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4277  (.I0(\edb_top_inst/n2945 ), .I1(\edb_top_inst/la0/data_out_shift_reg[20] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4277 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4278  (.I0(\edb_top_inst/la0/la_trig_mask[20] ), 
            .I1(\edb_top_inst/la0/la_run_trig ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2946 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4278 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__4279  (.I0(\edb_top_inst/n2946 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[20] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2947 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4279 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4280  (.I0(\edb_top_inst/n2947 ), .I1(\edb_top_inst/la0/data_out_shift_reg[21] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4280 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4281  (.I0(\edb_top_inst/la0/la_trig_mask[21] ), 
            .I1(\edb_top_inst/la0/la_run_trig_imdt ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2948 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4281 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__4282  (.I0(\edb_top_inst/la0/data_from_biu[21] ), 
            .I1(\edb_top_inst/n2948 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2949 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4282 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4283  (.I0(\edb_top_inst/n2949 ), .I1(\edb_top_inst/la0/data_out_shift_reg[22] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2445 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4283 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4284  (.I0(\edb_top_inst/la0/la_stop_trig ), 
            .I1(\edb_top_inst/n2901 ), .I2(\edb_top_inst/n2852 ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2950 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4284 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4285  (.I0(\edb_top_inst/la0/la_trig_mask[22] ), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/la0/data_from_biu[22] ), 
            .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2951 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4285 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__4286  (.I0(\edb_top_inst/n2950 ), .I1(\edb_top_inst/n2951 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[23] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4286 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4287  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[23] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2952 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4287 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4288  (.I0(\edb_top_inst/la0/data_from_biu[23] ), 
            .I1(\edb_top_inst/n2952 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2953 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4288 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4289  (.I0(\edb_top_inst/n2953 ), .I1(\edb_top_inst/la0/data_out_shift_reg[24] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4289 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4290  (.I0(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[24] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2954 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4290 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4291  (.I0(\edb_top_inst/n2954 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[24] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2955 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4291 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4292  (.I0(\edb_top_inst/n2955 ), .I1(\edb_top_inst/la0/data_out_shift_reg[25] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4292 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4293  (.I0(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[25] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2956 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4293 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4294  (.I0(\edb_top_inst/n2956 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[25] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2957 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4294 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4295  (.I0(\edb_top_inst/n2957 ), .I1(\edb_top_inst/la0/data_out_shift_reg[26] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4295 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4296  (.I0(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[26] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2958 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4296 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4297  (.I0(\edb_top_inst/n2958 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[26] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2959 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4297 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4298  (.I0(\edb_top_inst/n2959 ), .I1(\edb_top_inst/la0/data_out_shift_reg[27] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4298 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4299  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[27] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2960 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4299 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4300  (.I0(\edb_top_inst/la0/data_from_biu[27] ), 
            .I1(\edb_top_inst/n2960 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2961 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4300 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4301  (.I0(\edb_top_inst/n2961 ), .I1(\edb_top_inst/la0/data_out_shift_reg[28] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4301 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4302  (.I0(\edb_top_inst/la0/la_trig_pos[5] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[28] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2962 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4302 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4303  (.I0(\edb_top_inst/la0/data_from_biu[28] ), 
            .I1(\edb_top_inst/n2962 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2963 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4303 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4304  (.I0(\edb_top_inst/n2963 ), .I1(\edb_top_inst/la0/data_out_shift_reg[29] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4304 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4305  (.I0(\edb_top_inst/la0/la_trig_pos[6] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[29] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2964 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4305 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4306  (.I0(\edb_top_inst/la0/data_from_biu[29] ), 
            .I1(\edb_top_inst/n2964 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2965 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4306 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4307  (.I0(\edb_top_inst/n2965 ), .I1(\edb_top_inst/la0/data_out_shift_reg[30] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4307 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4308  (.I0(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[30] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2966 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4308 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4309  (.I0(\edb_top_inst/n2966 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[30] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2967 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4309 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4310  (.I0(\edb_top_inst/n2967 ), .I1(\edb_top_inst/la0/data_out_shift_reg[31] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4310 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4311  (.I0(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[31] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2968 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4311 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4312  (.I0(\edb_top_inst/la0/data_from_biu[31] ), 
            .I1(\edb_top_inst/n2968 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2969 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4312 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4313  (.I0(\edb_top_inst/n2969 ), .I1(\edb_top_inst/la0/data_out_shift_reg[32] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4313 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4314  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/n2901 ), .I2(\edb_top_inst/n2852 ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2970 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4314 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4315  (.I0(\edb_top_inst/la0/la_trig_mask[32] ), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/la0/data_from_biu[32] ), 
            .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2971 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4315 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__4316  (.I0(\edb_top_inst/n2970 ), .I1(\edb_top_inst/n2971 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[33] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4316 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4317  (.I0(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I1(\edb_top_inst/n2901 ), .I2(\edb_top_inst/n2852 ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2972 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4317 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4318  (.I0(\edb_top_inst/la0/la_trig_mask[33] ), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/la0/data_from_biu[33] ), 
            .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2973 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4318 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__4319  (.I0(\edb_top_inst/n2972 ), .I1(\edb_top_inst/n2973 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[34] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4319 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4320  (.I0(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[34] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2974 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4320 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4321  (.I0(\edb_top_inst/la0/data_from_biu[34] ), 
            .I1(\edb_top_inst/n2974 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2975 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4321 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4322  (.I0(\edb_top_inst/n2975 ), .I1(\edb_top_inst/la0/data_out_shift_reg[35] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4322 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4323  (.I0(\edb_top_inst/la0/la_trig_pos[12] ), 
            .I1(\edb_top_inst/n2901 ), .I2(\edb_top_inst/n2852 ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2976 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4323 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4324  (.I0(\edb_top_inst/la0/la_trig_mask[35] ), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/la0/data_from_biu[35] ), 
            .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2977 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4324 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__4325  (.I0(\edb_top_inst/n2976 ), .I1(\edb_top_inst/n2977 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[36] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4325 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4326  (.I0(\edb_top_inst/la0/la_trig_pos[13] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[36] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2978 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4326 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4327  (.I0(\edb_top_inst/la0/data_from_biu[36] ), 
            .I1(\edb_top_inst/n2978 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2979 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4327 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4328  (.I0(\edb_top_inst/n2979 ), .I1(\edb_top_inst/la0/data_out_shift_reg[37] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4328 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4329  (.I0(\edb_top_inst/la0/la_trig_pos[14] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[37] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2980 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4329 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4330  (.I0(\edb_top_inst/n2980 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[37] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2981 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4330 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4331  (.I0(\edb_top_inst/n2981 ), .I1(\edb_top_inst/la0/data_out_shift_reg[38] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4331 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4332  (.I0(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[38] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2982 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4332 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4333  (.I0(\edb_top_inst/n2982 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[38] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2983 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4333 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4334  (.I0(\edb_top_inst/n2983 ), .I1(\edb_top_inst/la0/data_out_shift_reg[39] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4334 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4335  (.I0(\edb_top_inst/la0/la_trig_pos[16] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[39] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2984 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4335 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4336  (.I0(\edb_top_inst/n2984 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[39] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2985 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4336 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4337  (.I0(\edb_top_inst/n2985 ), .I1(\edb_top_inst/la0/data_out_shift_reg[40] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4337 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4338  (.I0(\edb_top_inst/la0/la_trig_mask[40] ), 
            .I1(\edb_top_inst/la0/la_trig_pattern[0] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2986 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4338 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__4339  (.I0(\edb_top_inst/la0/data_from_biu[40] ), 
            .I1(\edb_top_inst/n2986 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2987 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4339 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4340  (.I0(\edb_top_inst/n2987 ), .I1(\edb_top_inst/la0/data_out_shift_reg[41] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4340 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4341  (.I0(\edb_top_inst/la0/la_trig_pattern[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[41] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2988 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4341 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4342  (.I0(\edb_top_inst/n2988 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[41] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2989 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4342 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4343  (.I0(\edb_top_inst/n2989 ), .I1(\edb_top_inst/la0/data_out_shift_reg[42] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2425 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4343 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4344  (.I0(\edb_top_inst/la0/la_capture_pattern[0] ), 
            .I1(\edb_top_inst/n2901 ), .I2(\edb_top_inst/n2852 ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2990 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4344 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4345  (.I0(\edb_top_inst/la0/la_trig_mask[42] ), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/la0/data_from_biu[42] ), 
            .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2991 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4345 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__4346  (.I0(\edb_top_inst/n2990 ), .I1(\edb_top_inst/n2991 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[43] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4346 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4347  (.I0(\edb_top_inst/la0/la_capture_pattern[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[43] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2992 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4347 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4348  (.I0(\edb_top_inst/n2855 ), .I1(\edb_top_inst/n2992 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[44] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2423 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf088, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4348 .LUTMASK = 16'hf088;
    EFX_LUT4 \edb_top_inst/LUT__4349  (.I0(\edb_top_inst/n2855 ), .I1(\edb_top_inst/n2853 ), 
            .O(\edb_top_inst/n2993 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4349 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4350  (.I0(\edb_top_inst/n2993 ), .I1(\edb_top_inst/la0/la_trig_mask[44] ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[45] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf088, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4350 .LUTMASK = 16'hf088;
    EFX_LUT4 \edb_top_inst/LUT__4351  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[45] ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2994 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4351 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4352  (.I0(\edb_top_inst/la0/data_out_shift_reg[46] ), 
            .I1(\edb_top_inst/n2994 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2421 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4352 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4353  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[46] ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2995 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4353 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4354  (.I0(\edb_top_inst/la0/data_out_shift_reg[47] ), 
            .I1(\edb_top_inst/n2995 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4354 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4355  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[47] ), .I2(\edb_top_inst/n2901 ), 
            .I3(\edb_top_inst/n2852 ), .O(\edb_top_inst/n2996 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4355 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4356  (.I0(\edb_top_inst/la0/data_out_shift_reg[48] ), 
            .I1(\edb_top_inst/n2996 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2419 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4356 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4357  (.I0(\edb_top_inst/n2993 ), .I1(\edb_top_inst/la0/la_trig_mask[48] ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[49] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf088, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4357 .LUTMASK = 16'hf088;
    EFX_LUT4 \edb_top_inst/LUT__4358  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[49] ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2997 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4358 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4359  (.I0(\edb_top_inst/la0/data_out_shift_reg[50] ), 
            .I1(\edb_top_inst/n2997 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2417 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4359 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4360  (.I0(\edb_top_inst/n2993 ), .I1(\edb_top_inst/la0/la_trig_mask[50] ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[51] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf088, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4360 .LUTMASK = 16'hf088;
    EFX_LUT4 \edb_top_inst/LUT__4361  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[51] ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2998 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4361 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4362  (.I0(\edb_top_inst/la0/data_out_shift_reg[52] ), 
            .I1(\edb_top_inst/n2998 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2415 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4362 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4363  (.I0(\edb_top_inst/n2993 ), .I1(\edb_top_inst/la0/la_trig_mask[52] ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[53] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf088, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4363 .LUTMASK = 16'hf088;
    EFX_LUT4 \edb_top_inst/LUT__4364  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[53] ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2999 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4364 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4365  (.I0(\edb_top_inst/la0/data_out_shift_reg[54] ), 
            .I1(\edb_top_inst/n2999 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2413 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4365 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4366  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[54] ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n3000 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4366 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4367  (.I0(\edb_top_inst/la0/data_out_shift_reg[55] ), 
            .I1(\edb_top_inst/n3000 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4367 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4368  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[55] ), .I2(\edb_top_inst/n2901 ), 
            .I3(\edb_top_inst/n2849 ), .O(\edb_top_inst/n3001 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4368 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4369  (.I0(\edb_top_inst/la0/data_out_shift_reg[56] ), 
            .I1(\edb_top_inst/n3001 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2411 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4369 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4370  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[56] ), .I2(\edb_top_inst/n2901 ), 
            .I3(\edb_top_inst/n2852 ), .O(\edb_top_inst/n3002 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4370 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4371  (.I0(\edb_top_inst/la0/data_out_shift_reg[57] ), 
            .I1(\edb_top_inst/n3002 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4371 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4372  (.I0(\edb_top_inst/n2993 ), .I1(\edb_top_inst/la0/la_trig_mask[57] ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[58] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2409 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf088, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4372 .LUTMASK = 16'hf088;
    EFX_LUT4 \edb_top_inst/LUT__4373  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[58] ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n3003 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4373 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4374  (.I0(\edb_top_inst/la0/data_out_shift_reg[59] ), 
            .I1(\edb_top_inst/n3003 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2408 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4374 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4375  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[59] ), .I2(\edb_top_inst/n2901 ), 
            .I3(\edb_top_inst/n2849 ), .O(\edb_top_inst/n3004 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4375 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4376  (.I0(\edb_top_inst/la0/data_out_shift_reg[60] ), 
            .I1(\edb_top_inst/n3004 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2407 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4376 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4377  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[60] ), .I2(\edb_top_inst/n2901 ), 
            .I3(\edb_top_inst/n2852 ), .O(\edb_top_inst/n3005 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4377 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4378  (.I0(\edb_top_inst/la0/data_out_shift_reg[61] ), 
            .I1(\edb_top_inst/n3005 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4378 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4379  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[61] ), .I2(\edb_top_inst/n2901 ), 
            .I3(\edb_top_inst/n2852 ), .O(\edb_top_inst/n3006 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4379 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4380  (.I0(\edb_top_inst/la0/data_out_shift_reg[62] ), 
            .I1(\edb_top_inst/n3006 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2405 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4380 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4381  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[62] ), .I2(\edb_top_inst/n2901 ), 
            .I3(\edb_top_inst/n2852 ), .O(\edb_top_inst/n3007 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4381 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4382  (.I0(\edb_top_inst/la0/data_out_shift_reg[63] ), 
            .I1(\edb_top_inst/n3007 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2404 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4382 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4383  (.I0(\edb_top_inst/la0/la_trig_mask[63] ), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/n2906 ), .O(\edb_top_inst/n3008 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4383 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4384  (.I0(\edb_top_inst/n2857 ), .I1(\edb_top_inst/n3008 ), 
            .I2(\edb_top_inst/n2901 ), .O(\edb_top_inst/la0/n2403 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4384 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4385  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/biu_ready ), .I2(jtag_inst2_UPDATE), .I3(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n3009 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f57, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4385 .LUTMASK = 16'h0f57;
    EFX_LUT4 \edb_top_inst/LUT__4386  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/n2839 ), .I2(\edb_top_inst/n2835 ), .I3(\edb_top_inst/n2811 ), 
            .O(\edb_top_inst/n3010 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4386 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4387  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/n3009 ), .I2(\edb_top_inst/n3010 ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n3011 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4387 .LUTMASK = 16'h00f8;
    EFX_LUT4 \edb_top_inst/LUT__4388  (.I0(\edb_top_inst/n2811 ), .I1(jtag_inst2_UPDATE), 
            .I2(\edb_top_inst/n2782 ), .I3(\edb_top_inst/n3011 ), .O(\edb_top_inst/la0/module_next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4388 .LUTMASK = 16'hff10;
    EFX_LUT4 \edb_top_inst/LUT__4389  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/n2823 ), 
            .I3(\edb_top_inst/n2828 ), .O(\edb_top_inst/n3012 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4389 .LUTMASK = 16'hb200;
    EFX_LUT4 \edb_top_inst/LUT__4390  (.I0(\edb_top_inst/n2830 ), .I1(\edb_top_inst/n3012 ), 
            .I2(\edb_top_inst/n2828 ), .I3(\edb_top_inst/n2835 ), .O(\edb_top_inst/n3013 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h30fa, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4390 .LUTMASK = 16'h30fa;
    EFX_LUT4 \edb_top_inst/LUT__4391  (.I0(\edb_top_inst/n2808 ), .I1(\edb_top_inst/n3013 ), 
            .I2(\edb_top_inst/n2811 ), .I3(jtag_inst2_UPDATE), .O(\edb_top_inst/la0/module_next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4391 .LUTMASK = 16'he0ee;
    EFX_LUT4 \edb_top_inst/LUT__4392  (.I0(\edb_top_inst/n2790 ), .I1(\edb_top_inst/n2835 ), 
            .I2(\edb_top_inst/n2782 ), .O(\edb_top_inst/n3014 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4392 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__4393  (.I0(\edb_top_inst/n2835 ), .I1(\edb_top_inst/n2829 ), 
            .I2(\edb_top_inst/n3014 ), .I3(jtag_inst2_UPDATE), .O(\edb_top_inst/la0/module_next_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4393 .LUTMASK = 16'h00f8;
    EFX_LUT4 \edb_top_inst/LUT__4394  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[1] ), .O(\edb_top_inst/la0/axi_crc_i/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4394 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4395  (.I0(\edb_top_inst/n2811 ), .I1(\edb_top_inst/n2782 ), 
            .I2(\edb_top_inst/la0/op_reg_en ), .I3(\edb_top_inst/n2834 ), 
            .O(\edb_top_inst/ceg_net221 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4395 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4396  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[2] ), .O(\edb_top_inst/la0/axi_crc_i/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4396 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4397  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[3] ), .O(\edb_top_inst/la0/axi_crc_i/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4397 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4398  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[4] ), .O(\edb_top_inst/la0/axi_crc_i/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4398 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4399  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[5] ), .O(\edb_top_inst/la0/axi_crc_i/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4399 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4400  (.I0(jtag_inst2_TDI), .I1(\edb_top_inst/la0/data_out_shift_reg[0] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/la0/crc_data_out[0] ), 
            .O(\edb_top_inst/n3015 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac53, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4400 .LUTMASK = 16'hac53;
    EFX_LUT4 \edb_top_inst/LUT__4401  (.I0(\edb_top_inst/n3015 ), .I1(\edb_top_inst/n2834 ), 
            .O(\edb_top_inst/n3016 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4401 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4402  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[6] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4402 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4403  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[7] ), .O(\edb_top_inst/la0/axi_crc_i/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4403 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4404  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[8] ), .O(\edb_top_inst/la0/axi_crc_i/n143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4404 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4405  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[9] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4405 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4406  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[10] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4406 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4407  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[11] ), .O(\edb_top_inst/la0/axi_crc_i/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4407 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4408  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[12] ), .O(\edb_top_inst/la0/axi_crc_i/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4408 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4409  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[13] ), .O(\edb_top_inst/la0/axi_crc_i/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4409 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4410  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[14] ), .O(\edb_top_inst/la0/axi_crc_i/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4410 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4411  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[15] ), .O(\edb_top_inst/la0/axi_crc_i/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4411 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4412  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[16] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4412 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4413  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[17] ), .O(\edb_top_inst/la0/axi_crc_i/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4413 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4414  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[18] ), .O(\edb_top_inst/la0/axi_crc_i/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4414 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4415  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[19] ), .O(\edb_top_inst/la0/axi_crc_i/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4415 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4416  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[20] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4416 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4417  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[21] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4417 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4418  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[22] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4418 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4419  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[23] ), .O(\edb_top_inst/la0/axi_crc_i/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4419 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4420  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[24] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4420 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4421  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[25] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4421 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4422  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[26] ), .O(\edb_top_inst/la0/axi_crc_i/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4422 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4423  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[27] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4423 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4424  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[28] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4424 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4425  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[29] ), .O(\edb_top_inst/la0/axi_crc_i/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4425 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4426  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[30] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4426 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4427  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[31] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4427 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4428  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .O(\edb_top_inst/la0/axi_crc_i/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4428 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4429  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/n2796 ), 
            .I3(\edb_top_inst/n2798 ), .O(\edb_top_inst/n3017 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4429 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4430  (.I0(\edb_top_inst/n3017 ), .I1(\edb_top_inst/n2870 ), 
            .O(\edb_top_inst/la0/n2766 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4430 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4431  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4431 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4432  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4432 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4433  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4433 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4434  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4434 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4435  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3018 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4435 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4436  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3019 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4436 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4437  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3020 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4437 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4438  (.I0(\edb_top_inst/n3019 ), .I1(\edb_top_inst/n3018 ), 
            .I2(\edb_top_inst/n3020 ), .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4438 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4439  (.I0(\edb_top_inst/n3017 ), .I1(\edb_top_inst/n2865 ), 
            .O(\edb_top_inst/la0/n3599 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4439 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4440  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4440 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4441  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4441 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4442  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4442 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4443  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4443 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4444  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3021 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4444 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4445  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3022 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4445 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4446  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3023 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4446 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4447  (.I0(\edb_top_inst/n3022 ), .I1(\edb_top_inst/n3021 ), 
            .I2(\edb_top_inst/n3023 ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4447 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4448  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/n3017 ), .I2(\edb_top_inst/edb_user_dr[71] ), 
            .I3(\edb_top_inst/edb_user_dr[72] ), .O(\edb_top_inst/la0/n4432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4448 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4449  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4449 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4450  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4450 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4451  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4451 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4452  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4452 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4453  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3024 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4453 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4454  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3025 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4454 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4455  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3026 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4455 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4456  (.I0(\edb_top_inst/n3025 ), .I1(\edb_top_inst/n3024 ), 
            .I2(\edb_top_inst/n3026 ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4456 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4457  (.I0(\edb_top_inst/n2796 ), .I1(\edb_top_inst/n2862 ), 
            .O(\edb_top_inst/la0/n5279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4457 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4458  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4458 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4459  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4459 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4460  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b22, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4460 .LUTMASK = 16'h2b22;
    EFX_LUT4 \edb_top_inst/LUT__4461  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/equal_9/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6ff6, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4461 .LUTMASK = 16'h6ff6;
    EFX_LUT4 \edb_top_inst/LUT__4462  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3027 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4462 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__4463  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/n3027 ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3028 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4463 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__4464  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n3029 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4464 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4465  (.I0(\edb_top_inst/n3027 ), .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n3029 ), .O(\edb_top_inst/n3030 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4c70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4465 .LUTMASK = 16'h4c70;
    EFX_LUT4 \edb_top_inst/LUT__4466  (.I0(\edb_top_inst/n3030 ), .I1(\edb_top_inst/n3028 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4466 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4467  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4467 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4468  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n9 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4468 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4469  (.I0(\edb_top_inst/n2864 ), .I1(\edb_top_inst/n2870 ), 
            .O(\edb_top_inst/la0/n6114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4469 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4470  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4470 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4471  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4471 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4472  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4472 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4473  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4473 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4474  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3031 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4474 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4475  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3032 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4475 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4476  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3033 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4476 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4477  (.I0(\edb_top_inst/n3032 ), .I1(\edb_top_inst/n3031 ), 
            .I2(\edb_top_inst/n3033 ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4477 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4478  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4478 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4479  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4479 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4480  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4480 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4481  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4481 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4482  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3034 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4482 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4483  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3035 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4483 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4484  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3036 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4484 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4485  (.I0(\edb_top_inst/n3035 ), .I1(\edb_top_inst/n3034 ), 
            .I2(\edb_top_inst/n3036 ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4485 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4486  (.I0(\edb_top_inst/n2796 ), .I1(\edb_top_inst/n2866 ), 
            .O(\edb_top_inst/la0/n7892 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4486 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4487  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4487 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4488  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4488 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4489  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/n3037 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4489 .LUTMASK = 16'h8eaf;
    EFX_LUT4 \edb_top_inst/LUT__4490  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), .O(\edb_top_inst/n3038 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4490 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4491  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3039 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4491 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4492  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), .O(\edb_top_inst/n3040 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4492 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4493  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), .O(\edb_top_inst/n3041 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4493 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4494  (.I0(\edb_top_inst/n3039 ), .I1(\edb_top_inst/n3038 ), 
            .I2(\edb_top_inst/n3040 ), .I3(\edb_top_inst/n3041 ), .O(\edb_top_inst/n3042 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4494 .LUTMASK = 16'hd000;
    EFX_LUT4 \edb_top_inst/LUT__4495  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n3043 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4495 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4496  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/n3044 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4496 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4497  (.I0(\edb_top_inst/n3043 ), .I1(\edb_top_inst/n3040 ), 
            .I2(\edb_top_inst/n3044 ), .O(\edb_top_inst/n3045 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4497 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4498  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), .O(\edb_top_inst/n3046 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4498 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4499  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n3047 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4499 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4500  (.I0(\edb_top_inst/n3042 ), .I1(\edb_top_inst/n3045 ), 
            .I2(\edb_top_inst/n3046 ), .I3(\edb_top_inst/n3047 ), .O(\edb_top_inst/n3048 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4500 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__4501  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] ), .O(\edb_top_inst/n3049 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4501 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4502  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/n3050 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4502 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4503  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/n3051 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4503 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4504  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] ), .I2(\edb_top_inst/n3050 ), 
            .I3(\edb_top_inst/n3051 ), .O(\edb_top_inst/n3052 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4504 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4505  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] ), .O(\edb_top_inst/n3053 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4505 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4506  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/n3054 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4506 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4507  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] ), .I2(\edb_top_inst/n3054 ), 
            .O(\edb_top_inst/n3055 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4507 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4508  (.I0(\edb_top_inst/n3053 ), .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I3(\edb_top_inst/n3055 ), .O(\edb_top_inst/n3056 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4508 .LUTMASK = 16'hb200;
    EFX_LUT4 \edb_top_inst/LUT__4509  (.I0(\edb_top_inst/n3048 ), .I1(\edb_top_inst/n3049 ), 
            .I2(\edb_top_inst/n3052 ), .I3(\edb_top_inst/n3056 ), .O(\edb_top_inst/n3057 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4509 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__4510  (.I0(\edb_top_inst/n3037 ), .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] ), .I3(\edb_top_inst/n3057 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4510 .LUTMASK = 16'h00b2;
    EFX_LUT4 \edb_top_inst/LUT__4511  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] ), .O(\edb_top_inst/n3058 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4511 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4512  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), .I2(\edb_top_inst/n3052 ), 
            .I3(\edb_top_inst/n3058 ), .O(\edb_top_inst/n3059 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4512 .LUTMASK = 16'hd000;
    EFX_LUT4 \edb_top_inst/LUT__4513  (.I0(\edb_top_inst/n3038 ), .I1(\edb_top_inst/n3039 ), 
            .I2(\edb_top_inst/n3043 ), .I3(\edb_top_inst/n3044 ), .O(\edb_top_inst/n3060 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4513 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4514  (.I0(\edb_top_inst/n3049 ), .I1(\edb_top_inst/n3047 ), 
            .I2(\edb_top_inst/n3046 ), .I3(\edb_top_inst/n3053 ), .O(\edb_top_inst/n3061 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4514 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4515  (.I0(\edb_top_inst/n3055 ), .I1(\edb_top_inst/n3060 ), 
            .I2(\edb_top_inst/n3061 ), .O(\edb_top_inst/n3062 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4515 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4516  (.I0(\edb_top_inst/n3059 ), .I1(\edb_top_inst/n3062 ), 
            .I2(\edb_top_inst/n3040 ), .I3(\edb_top_inst/n3041 ), .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/equal_9/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4516 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__4517  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] ), 
            .O(\edb_top_inst/n3063 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4517 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4518  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] ), 
            .O(\edb_top_inst/n3064 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4518 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4519  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] ), 
            .O(\edb_top_inst/n3065 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4519 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4520  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] ), 
            .O(\edb_top_inst/n3066 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4520 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4521  (.I0(\edb_top_inst/n3063 ), .I1(\edb_top_inst/n3064 ), 
            .I2(\edb_top_inst/n3065 ), .I3(\edb_top_inst/n3066 ), .O(\edb_top_inst/n3067 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4521 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4522  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .O(\edb_top_inst/n3068 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4522 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4523  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .O(\edb_top_inst/n3069 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4523 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4524  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .O(\edb_top_inst/n3070 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4524 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4525  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .O(\edb_top_inst/n3071 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4525 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4526  (.I0(\edb_top_inst/n3068 ), .I1(\edb_top_inst/n3069 ), 
            .I2(\edb_top_inst/n3070 ), .I3(\edb_top_inst/n3071 ), .O(\edb_top_inst/n3072 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4526 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4527  (.I0(\edb_top_inst/n3067 ), .I1(\edb_top_inst/n3072 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/n3073 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4527 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__4528  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .I3(\edb_top_inst/n3073 ), .O(\edb_top_inst/n3074 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc513, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4528 .LUTMASK = 16'hc513;
    EFX_LUT4 \edb_top_inst/LUT__4529  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n3075 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4529 .LUTMASK = 16'hccca;
    EFX_LUT4 \edb_top_inst/LUT__4530  (.I0(\edb_top_inst/n3075 ), .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/n3074 ), .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4530 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4531  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n71 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4531 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4532  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4532 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4533  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4533 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4534  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4534 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4535  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4535 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4536  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4536 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4537  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4537 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4538  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4538 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4539  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4539 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4540  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4540 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4541  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4541 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4542  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4542 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4543  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4543 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4544  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4544 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4545  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4545 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4546  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4546 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4547  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4547 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4548  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4548 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4549  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4549 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4550  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4550 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4551  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4551 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4552  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4552 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4553  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4553 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4554  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n29 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4554 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4555  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4555 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4556  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4556 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4557  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4557 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4558  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4558 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4559  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4559 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4560  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4560 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4561  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4561 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4562  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4562 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4563  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4563 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4564  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4564 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4565  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3076 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4565 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4566  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3077 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4566 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4567  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3078 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4567 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4568  (.I0(\edb_top_inst/n3077 ), .I1(\edb_top_inst/n3076 ), 
            .I2(\edb_top_inst/n3078 ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4568 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4569  (.I0(\edb_top_inst/n2869 ), .I1(\edb_top_inst/n2870 ), 
            .O(\edb_top_inst/la0/n9630 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4569 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4570  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4570 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4571  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4571 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4572  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), .O(\edb_top_inst/n3079 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4572 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4573  (.I0(\edb_top_inst/n3079 ), .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] ), .O(\edb_top_inst/n3080 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4573 .LUTMASK = 16'h7171;
    EFX_LUT4 \edb_top_inst/LUT__4574  (.I0(\edb_top_inst/n3080 ), .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] ), .O(\edb_top_inst/n3081 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4574 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4575  (.I0(\edb_top_inst/n3081 ), .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] ), .O(\edb_top_inst/n3082 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4575 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4576  (.I0(\edb_top_inst/n3082 ), .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] ), .O(\edb_top_inst/n3083 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4576 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4577  (.I0(\edb_top_inst/n3083 ), .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] ), .O(\edb_top_inst/n3084 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4577 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4578  (.I0(\edb_top_inst/n3084 ), .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] ), .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4578 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4579  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n3085 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4579 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4580  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/n3086 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4580 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4581  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3087 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4581 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4582  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n3088 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4582 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4583  (.I0(\edb_top_inst/n3085 ), .I1(\edb_top_inst/n3086 ), 
            .I2(\edb_top_inst/n3087 ), .I3(\edb_top_inst/n3088 ), .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/equal_9/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4583 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__4584  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n3089 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4584 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4585  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n3090 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4585 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4586  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .O(\edb_top_inst/n3091 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4586 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4587  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n3092 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4587 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4588  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n3093 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4588 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4589  (.I0(\edb_top_inst/n3090 ), .I1(\edb_top_inst/n3091 ), 
            .I2(\edb_top_inst/n3092 ), .I3(\edb_top_inst/n3093 ), .O(\edb_top_inst/n3094 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4589 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4590  (.I0(\edb_top_inst/n3089 ), .I1(\edb_top_inst/n3094 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3095 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4590 .LUTMASK = 16'h5c3f;
    EFX_LUT4 \edb_top_inst/LUT__4591  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n3096 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4591 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__4592  (.I0(\edb_top_inst/n3096 ), .I1(\edb_top_inst/n3095 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4592 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4593  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4593 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4594  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4594 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4595  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4595 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4596  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4596 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4597  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4597 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4598  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4598 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4599  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4599 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4600  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4600 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4601  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4601 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4602  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4602 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4603  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4603 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4604  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4604 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4605  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4605 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4606  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4606 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4607  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4607 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4608  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4608 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4609  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), .O(\edb_top_inst/n3097 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4609 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4610  (.I0(\edb_top_inst/n3097 ), .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] ), .O(\edb_top_inst/n3098 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4610 .LUTMASK = 16'h7171;
    EFX_LUT4 \edb_top_inst/LUT__4611  (.I0(\edb_top_inst/n3098 ), .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] ), .O(\edb_top_inst/n3099 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4611 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4612  (.I0(\edb_top_inst/n3099 ), .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] ), .O(\edb_top_inst/n3100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4612 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4613  (.I0(\edb_top_inst/n3100 ), .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] ), .O(\edb_top_inst/n3101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4613 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4614  (.I0(\edb_top_inst/n3101 ), .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] ), .O(\edb_top_inst/n3102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4614 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4615  (.I0(\edb_top_inst/n3102 ), .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] ), .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4615 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4616  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n3103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4616 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4617  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/n3104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4617 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4618  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4618 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4619  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n3106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4619 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4620  (.I0(\edb_top_inst/n3103 ), .I1(\edb_top_inst/n3104 ), 
            .I2(\edb_top_inst/n3105 ), .I3(\edb_top_inst/n3106 ), .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/equal_9/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4620 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__4621  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n3107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4621 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4622  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n3108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4622 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4623  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .O(\edb_top_inst/n3109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4623 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4624  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n3110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4624 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4625  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n3111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4625 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4626  (.I0(\edb_top_inst/n3108 ), .I1(\edb_top_inst/n3109 ), 
            .I2(\edb_top_inst/n3110 ), .I3(\edb_top_inst/n3111 ), .O(\edb_top_inst/n3112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4626 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4627  (.I0(\edb_top_inst/n3107 ), .I1(\edb_top_inst/n3112 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4627 .LUTMASK = 16'h5c3f;
    EFX_LUT4 \edb_top_inst/LUT__4628  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n3114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4628 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__4629  (.I0(\edb_top_inst/n3114 ), .I1(\edb_top_inst/n3113 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4629 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4630  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4630 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4631  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4631 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4632  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4632 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4633  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4633 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4634  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4634 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4635  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4635 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4636  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4636 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4637  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4637 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4638  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4638 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4639  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4639 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4640  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4640 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4641  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4641 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4642  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4642 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4643  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4643 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4644  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4644 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4645  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4645 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4646  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4646 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4647  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4647 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4648  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4648 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4649  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4649 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4650  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4650 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4651  (.I0(\edb_top_inst/n3116 ), .I1(\edb_top_inst/n3115 ), 
            .I2(\edb_top_inst/n3117 ), .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4651 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4652  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4652 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4653  (.I0(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4653 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4654  (.I0(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4654 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4655  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4655 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4656  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4656 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4657  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4657 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4658  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4658 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4659  (.I0(\edb_top_inst/n3119 ), .I1(\edb_top_inst/n3118 ), 
            .I2(\edb_top_inst/n3120 ), .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4659 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4660  (.I0(\edb_top_inst/la0/la_trig_mask[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[0] ), .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4660 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4661  (.I0(\edb_top_inst/la0/la_trig_mask[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4661 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4662  (.I0(\edb_top_inst/la0/la_trig_mask[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4662 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4663  (.I0(\edb_top_inst/la0/la_trig_mask[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[4] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4663 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4664  (.I0(\edb_top_inst/n3121 ), .I1(\edb_top_inst/n3122 ), 
            .I2(\edb_top_inst/n3123 ), .I3(\edb_top_inst/n3124 ), .O(\edb_top_inst/n3125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4664 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4665  (.I0(\edb_top_inst/la0/la_trig_mask[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4665 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4666  (.I0(\edb_top_inst/la0/la_trig_mask[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[6] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4666 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4667  (.I0(\edb_top_inst/n3125 ), .I1(\edb_top_inst/n3126 ), 
            .I2(\edb_top_inst/n3127 ), .O(\edb_top_inst/n3128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4667 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4668  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[11] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[4] ), .O(\edb_top_inst/n3129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4668 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4669  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[2] ), .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[0] ), .O(\edb_top_inst/n3130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4669 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4670  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[5] ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[3] ), .O(\edb_top_inst/n3131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4670 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4671  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[8] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[1] ), .O(\edb_top_inst/n3132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4671 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4672  (.I0(\edb_top_inst/n3129 ), .I1(\edb_top_inst/n3130 ), 
            .I2(\edb_top_inst/n3131 ), .I3(\edb_top_inst/n3132 ), .O(\edb_top_inst/n3133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4672 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4673  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[9] ), .O(\edb_top_inst/n3134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4673 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4674  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[10] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[6] ), .O(\edb_top_inst/n3135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4674 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4675  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[7] ), .I2(\edb_top_inst/n3134 ), 
            .I3(\edb_top_inst/n3135 ), .O(\edb_top_inst/n3136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4675 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__4676  (.I0(\edb_top_inst/n3133 ), .I1(\edb_top_inst/n3136 ), 
            .I2(\edb_top_inst/n3128 ), .I3(\edb_top_inst/la0/la_trig_pattern[0] ), 
            .O(\edb_top_inst/n3137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4676 .LUTMASK = 16'h7077;
    EFX_LUT4 \edb_top_inst/LUT__4677  (.I0(\edb_top_inst/n3128 ), .I1(\edb_top_inst/la0/la_trig_pattern[1] ), 
            .I2(\edb_top_inst/n3137 ), .O(\edb_top_inst/la0/trigger_tu/n89 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc1c1, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4677 .LUTMASK = 16'hc1c1;
    EFX_LUT4 \edb_top_inst/LUT__4678  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[1] ), .I2(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n3138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4678 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4679  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/la0/la_trig_pos[6] ), 
            .O(\edb_top_inst/n3139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4679 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4680  (.I0(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[8] ), .I2(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[10] ), .O(\edb_top_inst/n3140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4680 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4681  (.I0(\edb_top_inst/n3138 ), .I1(\edb_top_inst/n3139 ), 
            .I2(\edb_top_inst/n3140 ), .O(\edb_top_inst/n3141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4681 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4682  (.I0(\edb_top_inst/la0/la_trig_pos[13] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[14] ), .I2(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[16] ), .O(\edb_top_inst/n3142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4682 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4683  (.I0(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[12] ), .I2(\edb_top_inst/n3141 ), 
            .I3(\edb_top_inst/n3142 ), .O(\edb_top_inst/n3143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4683 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4684  (.I0(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_p2 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n3144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4684 .LUTMASK = 16'h0e0e;
    EFX_LUT4 \edb_top_inst/LUT__4685  (.I0(\edb_top_inst/n3144 ), .I1(\edb_top_inst/n3143 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n3145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4685 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4686  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[10] ), .O(\edb_top_inst/n3146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4686 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4687  (.I0(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[8] ), .I2(\edb_top_inst/n3138 ), 
            .I3(\edb_top_inst/n3139 ), .O(\edb_top_inst/n3147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4687 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4688  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/n3146 ), .I2(\edb_top_inst/n3147 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .O(\edb_top_inst/n3148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4688 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__4689  (.I0(\edb_top_inst/la0/la_trig_pos[12] ), 
            .I1(\edb_top_inst/n3141 ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[11] ), .O(\edb_top_inst/n3149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4689 .LUTMASK = 16'heb7e;
    EFX_LUT4 \edb_top_inst/LUT__4690  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n3150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4690 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4691  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[1] ), .O(\edb_top_inst/n3151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4691 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4692  (.I0(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I1(\edb_top_inst/n3150 ), .I2(\edb_top_inst/n3151 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .O(\edb_top_inst/n3152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4692 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__4693  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .I2(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .O(\edb_top_inst/n3153 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4693 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__4694  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[6] ), .O(\edb_top_inst/n3154 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4694 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4695  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/n3138 ), 
            .I3(\edb_top_inst/n3154 ), .O(\edb_top_inst/n3155 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4695 .LUTMASK = 16'hef10;
    EFX_LUT4 \edb_top_inst/LUT__4696  (.I0(\edb_top_inst/n3152 ), .I1(\edb_top_inst/n3153 ), 
            .I2(\edb_top_inst/n3155 ), .I3(\edb_top_inst/n3142 ), .O(\edb_top_inst/n3156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4696 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4697  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[8] ), .O(\edb_top_inst/n3157 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4697 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4698  (.I0(\edb_top_inst/n3138 ), .I1(\edb_top_inst/n3139 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[7] ), .I3(\edb_top_inst/n3157 ), 
            .O(\edb_top_inst/n3158 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4698 .LUTMASK = 16'h8700;
    EFX_LUT4 \edb_top_inst/LUT__4699  (.I0(\edb_top_inst/n3138 ), .I1(\edb_top_inst/n3139 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[7] ), .I3(\edb_top_inst/n3157 ), 
            .O(\edb_top_inst/n3159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8ff7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4699 .LUTMASK = 16'h8ff7;
    EFX_LUT4 \edb_top_inst/LUT__4700  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .O(\edb_top_inst/n3160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4700 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4701  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/n3160 ), .I2(\edb_top_inst/n3138 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .O(\edb_top_inst/n3161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4701 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__4702  (.I0(\edb_top_inst/n3159 ), .I1(\edb_top_inst/n3158 ), 
            .I2(\edb_top_inst/n3161 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .O(\edb_top_inst/n3162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4702 .LUTMASK = 16'h050c;
    EFX_LUT4 \edb_top_inst/LUT__4703  (.I0(\edb_top_inst/n3148 ), .I1(\edb_top_inst/n3149 ), 
            .I2(\edb_top_inst/n3156 ), .I3(\edb_top_inst/n3162 ), .O(\edb_top_inst/n3163 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4703 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4704  (.I0(\edb_top_inst/n3163 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/n3145 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n3164 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4704 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__4705  (.I0(\edb_top_inst/la0/tu_trigger ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n3165 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4705 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4706  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n3166 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4706 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4707  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_trig_pos[8] ), 
            .O(\edb_top_inst/n3167 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf40b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4707 .LUTMASK = 16'hf40b;
    EFX_LUT4 \edb_top_inst/LUT__4708  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n3168 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4708 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4709  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n3169 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4709 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4710  (.I0(\edb_top_inst/n3168 ), .I1(\edb_top_inst/n3169 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_trig_pos[14] ), 
            .O(\edb_top_inst/n3170 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf807, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4710 .LUTMASK = 16'hf807;
    EFX_LUT4 \edb_top_inst/LUT__4711  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4711 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4712  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n3172 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4712 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4713  (.I0(\edb_top_inst/n3168 ), .I1(\edb_top_inst/n3171 ), 
            .I2(\edb_top_inst/n3172 ), .O(\edb_top_inst/n3173 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4713 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4714  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/la0/la_window_depth[4] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[16] ), .O(\edb_top_inst/n3174 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4714 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__4715  (.I0(\edb_top_inst/n3174 ), .I1(\edb_top_inst/n3173 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[6] ), .I3(\edb_top_inst/n3170 ), 
            .O(\edb_top_inst/n3175 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4715 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__4716  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n3176 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6ffc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4716 .LUTMASK = 16'h6ffc;
    EFX_LUT4 \edb_top_inst/LUT__4717  (.I0(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/n3176 ), 
            .I3(\edb_top_inst/n3171 ), .O(\edb_top_inst/n3177 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4717 .LUTMASK = 16'hf077;
    EFX_LUT4 \edb_top_inst/LUT__4718  (.I0(\edb_top_inst/n3177 ), .I1(\edb_top_inst/n3175 ), 
            .I2(\edb_top_inst/n3167 ), .O(\edb_top_inst/n3178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4718 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4719  (.I0(\edb_top_inst/la0/la_stop_trig ), 
            .I1(\edb_top_inst/n3165 ), .O(\edb_top_inst/n3179 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4719 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4720  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4720 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4721  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[13] ), .I2(\edb_top_inst/n3180 ), 
            .O(\edb_top_inst/n3181 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4721 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4722  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n3182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4722 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4723  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/n3171 ), .I3(\edb_top_inst/la0/la_trig_pos[4] ), 
            .O(\edb_top_inst/n3183 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4fb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4723 .LUTMASK = 16'h4fb0;
    EFX_LUT4 \edb_top_inst/LUT__4724  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[13] ), .O(\edb_top_inst/n3184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f82, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4724 .LUTMASK = 16'h7f82;
    EFX_LUT4 \edb_top_inst/LUT__4725  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n3185 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4725 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4726  (.I0(\edb_top_inst/n3185 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/n3184 ), .I3(\edb_top_inst/la0/la_trig_pos[9] ), 
            .O(\edb_top_inst/n3186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4726 .LUTMASK = 16'h0c0b;
    EFX_LUT4 \edb_top_inst/LUT__4727  (.I0(\edb_top_inst/n3186 ), .I1(\edb_top_inst/n3181 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/n3183 ), 
            .O(\edb_top_inst/n3187 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4727 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4728  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/n3169 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_trig_pos[12] ), 
            .O(\edb_top_inst/n3188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bf4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4728 .LUTMASK = 16'h0bf4;
    EFX_LUT4 \edb_top_inst/LUT__4729  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/n3172 ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[2] ), .O(\edb_top_inst/n3189 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4729 .LUTMASK = 16'h40bf;
    EFX_LUT4 \edb_top_inst/LUT__4730  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3190 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4730 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4731  (.I0(\edb_top_inst/n3189 ), .I1(\edb_top_inst/n3190 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[1] ), .O(\edb_top_inst/n3191 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7e7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4731 .LUTMASK = 16'he7e7;
    EFX_LUT4 \edb_top_inst/LUT__4732  (.I0(\edb_top_inst/n3169 ), .I1(\edb_top_inst/la0/la_window_depth[4] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[15] ), .I3(\edb_top_inst/la0/la_trig_pos[11] ), 
            .O(\edb_top_inst/n3192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3dfe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4732 .LUTMASK = 16'h3dfe;
    EFX_LUT4 \edb_top_inst/LUT__4733  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[0] ), .I3(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3193 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4733 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__4734  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4734 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4735  (.I0(\edb_top_inst/n3168 ), .I1(\edb_top_inst/n3194 ), 
            .I2(\edb_top_inst/n3171 ), .O(\edb_top_inst/n3195 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4735 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4736  (.I0(\edb_top_inst/n3192 ), .I1(\edb_top_inst/n3193 ), 
            .I2(\edb_top_inst/n3195 ), .I3(\edb_top_inst/la0/la_trig_pos[10] ), 
            .O(\edb_top_inst/n3196 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4736 .LUTMASK = 16'h1001;
    EFX_LUT4 \edb_top_inst/LUT__4737  (.I0(\edb_top_inst/n3188 ), .I1(\edb_top_inst/n3191 ), 
            .I2(\edb_top_inst/n3187 ), .I3(\edb_top_inst/n3196 ), .O(\edb_top_inst/n3197 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4737 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4738  (.I0(\edb_top_inst/n3165 ), .I1(\edb_top_inst/n3178 ), 
            .I2(\edb_top_inst/n3197 ), .I3(\edb_top_inst/n3179 ), .O(\edb_top_inst/n3198 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4738 .LUTMASK = 16'h00bf;
    EFX_LUT4 \edb_top_inst/LUT__4739  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/n3198 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/n3164 ), .O(\edb_top_inst/n3199 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4739 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__4740  (.I0(\edb_top_inst/n3194 ), .I1(\edb_top_inst/n3168 ), 
            .O(\edb_top_inst/n3200 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4740 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4741  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n3201 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4741 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4742  (.I0(\edb_top_inst/n3201 ), .I1(\edb_top_inst/n3166 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3202 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4742 .LUTMASK = 16'h0a03;
    EFX_LUT4 \edb_top_inst/LUT__4743  (.I0(\edb_top_inst/n3200 ), .I1(\edb_top_inst/n3202 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .O(\edb_top_inst/n3203 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4743 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__4744  (.I0(\edb_top_inst/n3172 ), .I1(\edb_top_inst/n3168 ), 
            .O(\edb_top_inst/n3204 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4744 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4745  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/n3172 ), 
            .O(\edb_top_inst/n3205 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4745 .LUTMASK = 16'h6060;
    EFX_LUT4 \edb_top_inst/LUT__4746  (.I0(\edb_top_inst/n3204 ), .I1(\edb_top_inst/n3205 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .O(\edb_top_inst/n3206 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4746 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__4747  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I3(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3207 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdcf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4747 .LUTMASK = 16'hbdcf;
    EFX_LUT4 \edb_top_inst/LUT__4748  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3208 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4748 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4749  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3209 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4749 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4750  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/n3209 ), 
            .O(\edb_top_inst/n3210 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4750 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4751  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/n3185 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .I3(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n3211 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4751 .LUTMASK = 16'h0c0b;
    EFX_LUT4 \edb_top_inst/LUT__4752  (.I0(\edb_top_inst/n3210 ), .I1(\edb_top_inst/n3211 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .O(\edb_top_inst/n3212 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1428, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4752 .LUTMASK = 16'h1428;
    EFX_LUT4 \edb_top_inst/LUT__4753  (.I0(\edb_top_inst/n3207 ), .I1(\edb_top_inst/n3208 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), .I3(\edb_top_inst/n3212 ), 
            .O(\edb_top_inst/n3213 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4753 .LUTMASK = 16'h1400;
    EFX_LUT4 \edb_top_inst/LUT__4754  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n3166 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n3214 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4754 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4755  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n3182 ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n3215 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4551, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4755 .LUTMASK = 16'h4551;
    EFX_LUT4 \edb_top_inst/LUT__4756  (.I0(\edb_top_inst/n3214 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), .I3(\edb_top_inst/n3215 ), 
            .O(\edb_top_inst/n3216 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4756 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__4757  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/n3171 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .O(\edb_top_inst/n3217 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4fb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4757 .LUTMASK = 16'h4fb0;
    EFX_LUT4 \edb_top_inst/LUT__4758  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/n3173 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), .I3(\edb_top_inst/n3217 ), 
            .O(\edb_top_inst/n3218 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3edf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4758 .LUTMASK = 16'h3edf;
    EFX_LUT4 \edb_top_inst/LUT__4759  (.I0(\edb_top_inst/n3216 ), .I1(\edb_top_inst/n3218 ), 
            .O(\edb_top_inst/n3219 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4759 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4760  (.I0(\edb_top_inst/n3203 ), .I1(\edb_top_inst/n3206 ), 
            .I2(\edb_top_inst/n3213 ), .I3(\edb_top_inst/n3219 ), .O(\edb_top_inst/n3220 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4760 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4761  (.I0(\edb_top_inst/n3168 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), .I3(\edb_top_inst/n3172 ), 
            .O(\edb_top_inst/n3221 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4761 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__4762  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
            .I3(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3222 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4762 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__4763  (.I0(\edb_top_inst/n3221 ), .I1(\edb_top_inst/n3222 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), .I3(\edb_top_inst/n3209 ), 
            .O(\edb_top_inst/n3223 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4763 .LUTMASK = 16'h0110;
    EFX_LUT4 \edb_top_inst/LUT__4764  (.I0(\edb_top_inst/n3214 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .O(\edb_top_inst/n3224 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4764 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4765  (.I0(\edb_top_inst/n3194 ), .I1(\edb_top_inst/n3171 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .O(\edb_top_inst/n3225 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4765 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__4766  (.I0(\edb_top_inst/n3201 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .O(\edb_top_inst/n3226 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf40b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4766 .LUTMASK = 16'hf40b;
    EFX_LUT4 \edb_top_inst/LUT__4767  (.I0(\edb_top_inst/n3168 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/n3171 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .O(\edb_top_inst/n3227 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4767 .LUTMASK = 16'h8f70;
    EFX_LUT4 \edb_top_inst/LUT__4768  (.I0(\edb_top_inst/n3225 ), .I1(\edb_top_inst/n3217 ), 
            .I2(\edb_top_inst/n3226 ), .I3(\edb_top_inst/n3227 ), .O(\edb_top_inst/n3228 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4768 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4769  (.I0(\edb_top_inst/n3169 ), .I1(\edb_top_inst/n3182 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3229 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4769 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4770  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n3185 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n3230 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4770 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4771  (.I0(\edb_top_inst/n3229 ), .I1(\edb_top_inst/n3230 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] ), 
            .O(\edb_top_inst/n3231 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1428, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4771 .LUTMASK = 16'h1428;
    EFX_LUT4 \edb_top_inst/LUT__4772  (.I0(\edb_top_inst/n3223 ), .I1(\edb_top_inst/n3224 ), 
            .I2(\edb_top_inst/n3228 ), .I3(\edb_top_inst/n3231 ), .O(\edb_top_inst/n3232 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4772 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4773  (.I0(\edb_top_inst/n3204 ), .I1(\edb_top_inst/n3205 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[3] ), .I3(\edb_top_inst/la0/la_trig_pos[2] ), 
            .O(\edb_top_inst/n3233 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4773 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__4774  (.I0(\edb_top_inst/n3200 ), .I1(\edb_top_inst/n3202 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[11] ), .I3(\edb_top_inst/la0/la_trig_pos[10] ), 
            .O(\edb_top_inst/n3234 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4774 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__4775  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/n3180 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[15] ), .O(\edb_top_inst/n3235 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ff4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4775 .LUTMASK = 16'h3ff4;
    EFX_LUT4 \edb_top_inst/LUT__4776  (.I0(\edb_top_inst/n3235 ), .I1(\edb_top_inst/n3230 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[9] ), .I3(\edb_top_inst/n3167 ), 
            .O(\edb_top_inst/n3236 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4776 .LUTMASK = 16'h1400;
    EFX_LUT4 \edb_top_inst/LUT__4777  (.I0(\edb_top_inst/n3233 ), .I1(\edb_top_inst/n3234 ), 
            .I2(\edb_top_inst/n3175 ), .I3(\edb_top_inst/n3236 ), .O(\edb_top_inst/n3237 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4777 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4778  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n3238 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4778 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4779  (.I0(\edb_top_inst/n3238 ), .I1(\edb_top_inst/la0/la_trig_pos[5] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[4] ), .I3(\edb_top_inst/n3210 ), 
            .O(\edb_top_inst/n3239 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4779 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__4780  (.I0(\edb_top_inst/n3185 ), .I1(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[1] ), .I3(\edb_top_inst/n3208 ), 
            .O(\edb_top_inst/n3240 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4780 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__4781  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n3169 ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3241 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4781 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4782  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/n3241 ), .I2(\edb_top_inst/la0/la_trig_pos[13] ), 
            .O(\edb_top_inst/n3242 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4782 .LUTMASK = 16'h1414;
    EFX_LUT4 \edb_top_inst/LUT__4783  (.I0(\edb_top_inst/n3239 ), .I1(\edb_top_inst/n3240 ), 
            .I2(\edb_top_inst/n3188 ), .I3(\edb_top_inst/n3242 ), .O(\edb_top_inst/n3243 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4783 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4784  (.I0(\edb_top_inst/n3232 ), .I1(\edb_top_inst/n3237 ), 
            .I2(\edb_top_inst/n3243 ), .O(\edb_top_inst/n3244 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4784 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4785  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[5] ), .I2(\edb_top_inst/la0/la_num_trigger[6] ), 
            .O(\edb_top_inst/n3245 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4785 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4786  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .I2(\edb_top_inst/la0/la_num_trigger[2] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[3] ), .O(\edb_top_inst/n3246 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4786 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4787  (.I0(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[8] ), .I2(\edb_top_inst/la0/la_num_trigger[9] ), 
            .O(\edb_top_inst/n3247 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4787 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4788  (.I0(\edb_top_inst/n3245 ), .I1(\edb_top_inst/n3246 ), 
            .I2(\edb_top_inst/n3247 ), .O(\edb_top_inst/n3248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4788 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4789  (.I0(\edb_top_inst/la0/la_num_trigger[11] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] ), .O(\edb_top_inst/n3249 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4789 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4790  (.I0(\edb_top_inst/la0/la_num_trigger[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), .I2(\edb_top_inst/n3248 ), 
            .I3(\edb_top_inst/n3249 ), .O(\edb_top_inst/n3250 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd6bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4790 .LUTMASK = 16'hd6bf;
    EFX_LUT4 \edb_top_inst/LUT__4791  (.I0(\edb_top_inst/n3249 ), .I1(\edb_top_inst/la0/la_num_trigger[10] ), 
            .I2(\edb_top_inst/la0/la_num_trigger[11] ), .I3(\edb_top_inst/la0/la_num_trigger[12] ), 
            .O(\edb_top_inst/n3251 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe45, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4791 .LUTMASK = 16'hfe45;
    EFX_LUT4 \edb_top_inst/LUT__4792  (.I0(\edb_top_inst/la0/la_num_trigger[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .O(\edb_top_inst/n3252 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4792 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4793  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .O(\edb_top_inst/n3253 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4793 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4794  (.I0(\edb_top_inst/la0/la_num_trigger[2] ), 
            .I1(\edb_top_inst/n3252 ), .I2(\edb_top_inst/n3253 ), .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .O(\edb_top_inst/n3254 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4794 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__4795  (.I0(\edb_top_inst/n3251 ), .I1(\edb_top_inst/n3254 ), 
            .O(\edb_top_inst/n3255 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4795 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4796  (.I0(\edb_top_inst/n3246 ), .I1(\edb_top_inst/n3245 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), .I3(\edb_top_inst/la0/la_num_trigger[7] ), 
            .O(\edb_top_inst/n3256 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h87f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4796 .LUTMASK = 16'h87f8;
    EFX_LUT4 \edb_top_inst/LUT__4797  (.I0(\edb_top_inst/la0/la_num_trigger[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .I2(\edb_top_inst/la0/la_num_trigger[9] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), .O(\edb_top_inst/n3257 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4797 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4798  (.I0(\edb_top_inst/la0/la_num_trigger[8] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[9] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .O(\edb_top_inst/n3258 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4798 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__4799  (.I0(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I1(\edb_top_inst/n3245 ), .I2(\edb_top_inst/n3246 ), .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .O(\edb_top_inst/n3259 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4799 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4800  (.I0(\edb_top_inst/n3258 ), .I1(\edb_top_inst/n3259 ), 
            .I2(\edb_top_inst/n3256 ), .I3(\edb_top_inst/n3257 ), .O(\edb_top_inst/n3260 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4800 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4801  (.I0(\edb_top_inst/la0/la_num_trigger[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), .O(\edb_top_inst/n3261 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4801 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4802  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/n3261 ), .I2(\edb_top_inst/n3246 ), .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .O(\edb_top_inst/n3262 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4802 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__4803  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[5] ), .I2(\edb_top_inst/n3246 ), 
            .I3(\edb_top_inst/la0/la_num_trigger[6] ), .O(\edb_top_inst/n3263 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4803 .LUTMASK = 16'hef10;
    EFX_LUT4 \edb_top_inst/LUT__4804  (.I0(\edb_top_inst/la0/la_num_trigger[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .O(\edb_top_inst/n3264 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4804 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4805  (.I0(\edb_top_inst/la0/la_num_trigger[13] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[14] ), .I2(\edb_top_inst/la0/la_num_trigger[15] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[16] ), .O(\edb_top_inst/n3265 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4805 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4806  (.I0(\edb_top_inst/n3264 ), .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .I2(\edb_top_inst/la0/la_num_trigger[0] ), .I3(\edb_top_inst/n3265 ), 
            .O(\edb_top_inst/n3266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4806 .LUTMASK = 16'h1800;
    EFX_LUT4 \edb_top_inst/LUT__4807  (.I0(\edb_top_inst/n3262 ), .I1(\edb_top_inst/n3263 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .I3(\edb_top_inst/n3266 ), 
            .O(\edb_top_inst/n3267 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4807 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__4808  (.I0(\edb_top_inst/n3250 ), .I1(\edb_top_inst/n3260 ), 
            .I2(\edb_top_inst/n3255 ), .I3(\edb_top_inst/n3267 ), .O(\edb_top_inst/n3268 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4808 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4809  (.I0(\edb_top_inst/n3268 ), .I1(\edb_top_inst/n3143 ), 
            .O(\edb_top_inst/n3269 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4809 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4810  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n3270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4810 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4811  (.I0(\edb_top_inst/n3244 ), .I1(\edb_top_inst/n3220 ), 
            .I2(\edb_top_inst/n3269 ), .I3(\edb_top_inst/n3270 ), .O(\edb_top_inst/n3271 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4811 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4812  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/n3165 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3272 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4812 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__4813  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .O(\edb_top_inst/n3273 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4813 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4814  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/n3232 ), .I2(\edb_top_inst/n3272 ), .I3(\edb_top_inst/n3273 ), 
            .O(\edb_top_inst/n3274 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4814 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__4815  (.I0(\edb_top_inst/n3163 ), .I1(\edb_top_inst/n3273 ), 
            .I2(\edb_top_inst/n3274 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n3275 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4815 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4816  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/n3271 ), .I2(\edb_top_inst/n3199 ), .I3(\edb_top_inst/n3275 ), 
            .O(\edb_top_inst/la0/la_biu_inst/next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h10ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4816 .LUTMASK = 16'h10ff;
    EFX_LUT4 \edb_top_inst/LUT__4817  (.I0(\edb_top_inst/n2825 ), .I1(\edb_top_inst/n2818 ), 
            .I2(\edb_top_inst/la0/biu_ready ), .O(\edb_top_inst/la0/la_biu_inst/n382 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4817 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4818  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), .O(\edb_top_inst/la0/la_biu_inst/n1315 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4818 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4819  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), .I2(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q ), 
            .I3(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), .O(\edb_top_inst/la0/la_biu_inst/next_fsm_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00be, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4819 .LUTMASK = 16'h00be;
    EFX_LUT4 \edb_top_inst/LUT__4820  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .I2(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .O(\edb_top_inst/ceg_net351 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4820 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4821  (.I0(\edb_top_inst/n3165 ), .I1(\edb_top_inst/n3178 ), 
            .I2(\edb_top_inst/n3197 ), .O(\edb_top_inst/n3276 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4821 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4822  (.I0(\edb_top_inst/n3268 ), .I1(\edb_top_inst/n3165 ), 
            .O(\edb_top_inst/n3277 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4822 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4823  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3278 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4823 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4824  (.I0(\edb_top_inst/n3232 ), .I1(\edb_top_inst/n3277 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I3(\edb_top_inst/n3278 ), 
            .O(\edb_top_inst/n3279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4824 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4825  (.I0(\edb_top_inst/n2903 ), .I1(\edb_top_inst/n3276 ), 
            .I2(\edb_top_inst/n3271 ), .I3(\edb_top_inst/n3279 ), .O(\edb_top_inst/la0/la_biu_inst/n1300 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4825 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__4826  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/n17781 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4826 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4827  (.I0(\edb_top_inst/n3244 ), .I1(\edb_top_inst/n3220 ), 
            .I2(\edb_top_inst/n3269 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .O(\edb_top_inst/n3280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4827 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__4828  (.I0(\edb_top_inst/n3179 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n3281 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4828 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4829  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n3282 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4829 .LUTMASK = 16'h0e00;
    EFX_LUT4 \edb_top_inst/LUT__4830  (.I0(\edb_top_inst/n3276 ), .I1(\edb_top_inst/n3277 ), 
            .I2(\edb_top_inst/n3281 ), .I3(\edb_top_inst/n3282 ), .O(\edb_top_inst/n3283 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4830 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__4831  (.I0(\edb_top_inst/n3232 ), .I1(\edb_top_inst/n2904 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3284 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4831 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__4832  (.I0(\edb_top_inst/n3165 ), .I1(\edb_top_inst/n3278 ), 
            .I2(\edb_top_inst/n3268 ), .O(\edb_top_inst/n3285 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4832 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4833  (.I0(\edb_top_inst/n3285 ), .I1(\edb_top_inst/n3284 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n3286 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4833 .LUTMASK = 16'h0a0c;
    EFX_LUT4 \edb_top_inst/LUT__4834  (.I0(\edb_top_inst/n3280 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/n3283 ), .I3(\edb_top_inst/n3286 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4834 .LUTMASK = 16'hff0b;
    EFX_LUT4 \edb_top_inst/LUT__4835  (.I0(\edb_top_inst/n3144 ), .I1(\edb_top_inst/n3143 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I3(\edb_top_inst/n3163 ), 
            .O(\edb_top_inst/n3287 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4835 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4836  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/n3165 ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3288 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4836 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__4837  (.I0(\edb_top_inst/n2904 ), .I1(\edb_top_inst/n3232 ), 
            .I2(\edb_top_inst/n3288 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .O(\edb_top_inst/n3289 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4837 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__4838  (.I0(\edb_top_inst/n3287 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I3(\edb_top_inst/n3289 ), 
            .O(\edb_top_inst/n3290 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4838 .LUTMASK = 16'hf100;
    EFX_LUT4 \edb_top_inst/LUT__4839  (.I0(\edb_top_inst/n3179 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/n3277 ), .I3(\edb_top_inst/n3276 ), .O(\edb_top_inst/n3291 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4839 .LUTMASK = 16'h1001;
    EFX_LUT4 \edb_top_inst/LUT__4840  (.I0(\edb_top_inst/n3143 ), .I1(\edb_top_inst/n3268 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .O(\edb_top_inst/n3292 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4840 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__4841  (.I0(\edb_top_inst/n3288 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n3293 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4841 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4842  (.I0(\edb_top_inst/n3244 ), .I1(\edb_top_inst/n3220 ), 
            .I2(\edb_top_inst/n3292 ), .I3(\edb_top_inst/n3293 ), .O(\edb_top_inst/n3294 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4842 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__4843  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/n3163 ), .I2(\edb_top_inst/n3273 ), .O(\edb_top_inst/n3295 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4843 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__4844  (.I0(\edb_top_inst/n3294 ), .I1(\edb_top_inst/n3291 ), 
            .I2(\edb_top_inst/n3290 ), .I3(\edb_top_inst/n3295 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4844 .LUTMASK = 16'hfff2;
    EFX_LUT4 \edb_top_inst/LUT__4845  (.I0(\edb_top_inst/la0/la_biu_inst/n382 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), .I2(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q ), 
            .O(\edb_top_inst/ceg_net348 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4845 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__4846  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), .O(\edb_top_inst/la0/la_biu_inst/next_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4846 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4847  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/n3165 ), .I2(\edb_top_inst/n2903 ), .O(\edb_top_inst/la0/la_biu_inst/n2053 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4847 .LUTMASK = 16'hbfbf;
    EFX_LUT4 \edb_top_inst/LUT__4848  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/la0/la_biu_inst/fifo_push )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05fc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4848 .LUTMASK = 16'h05fc;
    EFX_LUT4 \edb_top_inst/LUT__4849  (.I0(\edb_top_inst/la0/la_biu_inst/n2053 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_push ), .O(\edb_top_inst/n3296 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4849 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4850  (.I0(\edb_top_inst/n3232 ), .I1(\edb_top_inst/n3296 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4850 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4851  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n3297 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4851 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4852  (.I0(\edb_top_inst/n3297 ), .I1(\edb_top_inst/la0/la_resetn ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_rstn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4852 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4853  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4853 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4854  (.I0(\edb_top_inst/n3296 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
            .O(\edb_top_inst/ceg_net355 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4854 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4855  (.I0(\edb_top_inst/n2909 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4855 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4856  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[15] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4856 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4857  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[16] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4857 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4858  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[17] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4858 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4859  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[18] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4859 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4860  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[19] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4860 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4861  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[20] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4861 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4862  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[21] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4862 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4863  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[22] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4863 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4864  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[23] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4864 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4865  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[24] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4865 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4866  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[25] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4866 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4867  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[26] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4867 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4868  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .O(\edb_top_inst/n3298 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4868 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4869  (.I0(\edb_top_inst/n3172 ), .I1(\edb_top_inst/n3298 ), 
            .I2(\edb_top_inst/n3215 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4869 .LUTMASK = 16'hf888;
    EFX_LUT4 \edb_top_inst/LUT__4870  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .I3(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3299 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4870 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__4871  (.I0(\edb_top_inst/n3172 ), .I1(\edb_top_inst/n3299 ), 
            .O(\edb_top_inst/n3300 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4871 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4872  (.I0(\edb_top_inst/n3180 ), .I1(\edb_top_inst/n3229 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] ), 
            .I3(\edb_top_inst/n3300 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4872 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4873  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n3301 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4873 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4874  (.I0(\edb_top_inst/n3168 ), .I1(\edb_top_inst/n3301 ), 
            .I2(\edb_top_inst/n3229 ), .O(\edb_top_inst/n3302 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4874 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4875  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3303 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4875 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4876  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .I2(\edb_top_inst/n3303 ), 
            .I3(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3304 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4876 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4877  (.I0(\edb_top_inst/n3304 ), .I1(\edb_top_inst/n3172 ), 
            .I2(\edb_top_inst/n3302 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4877 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4878  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3305 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4878 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4879  (.I0(\edb_top_inst/n3305 ), .I1(\edb_top_inst/n3303 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3306 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4879 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4880  (.I0(\edb_top_inst/n3306 ), .I1(\edb_top_inst/n3172 ), 
            .O(\edb_top_inst/n3307 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4880 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4881  (.I0(\edb_top_inst/n3301 ), .I1(\edb_top_inst/n3229 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] ), 
            .I3(\edb_top_inst/n3307 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4881 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4882  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3308 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b04, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4882 .LUTMASK = 16'h0b04;
    EFX_LUT4 \edb_top_inst/LUT__4883  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3309 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4883 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4884  (.I0(\edb_top_inst/n3309 ), .I1(\edb_top_inst/n3305 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3310 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4884 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4885  (.I0(\edb_top_inst/n3310 ), .I1(\edb_top_inst/n3298 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3311 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4885 .LUTMASK = 16'hc500;
    EFX_LUT4 \edb_top_inst/LUT__4886  (.I0(\edb_top_inst/n3308 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] ), 
            .I2(\edb_top_inst/n3311 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4886 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4887  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3312 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4887 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4888  (.I0(\edb_top_inst/n3312 ), .I1(\edb_top_inst/n3309 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3313 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4888 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4889  (.I0(\edb_top_inst/n3299 ), .I1(\edb_top_inst/n3313 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3314 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4889 .LUTMASK = 16'ha300;
    EFX_LUT4 \edb_top_inst/LUT__4890  (.I0(\edb_top_inst/n3238 ), .I1(\edb_top_inst/n3308 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] ), 
            .I3(\edb_top_inst/n3314 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4890 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4891  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .I3(\edb_top_inst/n3308 ), .O(\edb_top_inst/n3315 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4891 .LUTMASK = 16'hd700;
    EFX_LUT4 \edb_top_inst/LUT__4892  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3316 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4892 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4893  (.I0(\edb_top_inst/n3316 ), .I1(\edb_top_inst/n3312 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3317 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4893 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4894  (.I0(\edb_top_inst/n3317 ), .I1(\edb_top_inst/n3304 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3318 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4894 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4895  (.I0(\edb_top_inst/n3315 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] ), 
            .I2(\edb_top_inst/n3318 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4895 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4896  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n3182 ), .I2(\edb_top_inst/n3308 ), .O(\edb_top_inst/n3319 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4896 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__4897  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3320 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4897 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4898  (.I0(\edb_top_inst/n3320 ), .I1(\edb_top_inst/n3316 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3321 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4898 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4899  (.I0(\edb_top_inst/n3321 ), .I1(\edb_top_inst/n3306 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3322 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4899 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4900  (.I0(\edb_top_inst/n3319 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] ), 
            .I2(\edb_top_inst/n3322 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4900 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4901  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3323 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4901 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4902  (.I0(\edb_top_inst/n3323 ), .I1(\edb_top_inst/n3320 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3324 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4902 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4903  (.I0(\edb_top_inst/n3324 ), .I1(\edb_top_inst/n3298 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3325 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf30a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4903 .LUTMASK = 16'hf30a;
    EFX_LUT4 \edb_top_inst/LUT__4904  (.I0(\edb_top_inst/n3310 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/n3325 ), 
            .O(\edb_top_inst/n3326 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4904 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4905  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/n3319 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] ), 
            .I3(\edb_top_inst/n3326 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4905 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4906  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3327 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4906 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4907  (.I0(\edb_top_inst/n3327 ), .I1(\edb_top_inst/n3323 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3328 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4907 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4908  (.I0(\edb_top_inst/n3328 ), .I1(\edb_top_inst/n3299 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3329 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf30a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4908 .LUTMASK = 16'hf30a;
    EFX_LUT4 \edb_top_inst/LUT__4909  (.I0(\edb_top_inst/n3313 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/n3329 ), 
            .O(\edb_top_inst/n3330 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4909 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4910  (.I0(\edb_top_inst/n3185 ), .I1(\edb_top_inst/n3319 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] ), 
            .I3(\edb_top_inst/n3330 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4910 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4911  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3331 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4911 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4912  (.I0(\edb_top_inst/n3331 ), .I1(\edb_top_inst/n3327 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3332 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4912 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4913  (.I0(\edb_top_inst/n3332 ), .I1(\edb_top_inst/n3317 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3333 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4913 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4914  (.I0(\edb_top_inst/n3304 ), .I1(\edb_top_inst/n3194 ), 
            .I2(\edb_top_inst/la0/la_window_depth[3] ), .I3(\edb_top_inst/n3333 ), 
            .O(\edb_top_inst/n3334 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4914 .LUTMASK = 16'h00bf;
    EFX_LUT4 \edb_top_inst/LUT__4915  (.I0(\edb_top_inst/n3201 ), .I1(\edb_top_inst/n3319 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] ), 
            .I3(\edb_top_inst/n3334 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4915 .LUTMASK = 16'h40ff;
    EFX_LUT4 \edb_top_inst/LUT__4916  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n3335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4916 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4917  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4917 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4918  (.I0(\edb_top_inst/n3336 ), .I1(\edb_top_inst/n3331 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3337 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4918 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4919  (.I0(\edb_top_inst/n3337 ), .I1(\edb_top_inst/n3321 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3338 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4919 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4920  (.I0(\edb_top_inst/n3306 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/n3194 ), .I3(\edb_top_inst/n3338 ), .O(\edb_top_inst/n3339 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4920 .LUTMASK = 16'h00bf;
    EFX_LUT4 \edb_top_inst/LUT__4921  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] ), 
            .I1(\edb_top_inst/n3308 ), .I2(\edb_top_inst/n3335 ), .I3(\edb_top_inst/n3339 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h80ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4921 .LUTMASK = 16'h80ff;
    EFX_LUT4 \edb_top_inst/LUT__4922  (.I0(\edb_top_inst/n3172 ), .I1(\edb_top_inst/n3298 ), 
            .I2(\edb_top_inst/n3215 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4922 .LUTMASK = 16'hf888;
    EFX_LUT4 \edb_top_inst/LUT__4923  (.I0(\edb_top_inst/n3180 ), .I1(\edb_top_inst/n3229 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] ), 
            .I3(\edb_top_inst/n3300 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4923 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4924  (.I0(\edb_top_inst/n3304 ), .I1(\edb_top_inst/n3172 ), 
            .I2(\edb_top_inst/n3302 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4924 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4925  (.I0(\edb_top_inst/n3301 ), .I1(\edb_top_inst/n3229 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] ), 
            .I3(\edb_top_inst/n3307 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4925 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4926  (.I0(\edb_top_inst/n3308 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] ), 
            .I2(\edb_top_inst/n3311 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4926 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4927  (.I0(\edb_top_inst/n3238 ), .I1(\edb_top_inst/n3308 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] ), 
            .I3(\edb_top_inst/n3314 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4927 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4928  (.I0(\edb_top_inst/n3315 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] ), 
            .I2(\edb_top_inst/n3318 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4928 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4929  (.I0(\edb_top_inst/n3319 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] ), 
            .I2(\edb_top_inst/n3322 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4929 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4930  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/n3319 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] ), 
            .I3(\edb_top_inst/n3326 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4930 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4931  (.I0(\edb_top_inst/n3185 ), .I1(\edb_top_inst/n3319 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] ), 
            .I3(\edb_top_inst/n3330 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4931 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4932  (.I0(\edb_top_inst/n3201 ), .I1(\edb_top_inst/n3319 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] ), 
            .I3(\edb_top_inst/n3334 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4932 .LUTMASK = 16'h40ff;
    EFX_LUT4 \edb_top_inst/LUT__4933  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] ), 
            .I1(\edb_top_inst/n3308 ), .I2(\edb_top_inst/n3335 ), .I3(\edb_top_inst/n3339 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h80ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4933 .LUTMASK = 16'h80ff;
    EFX_LUT4 \edb_top_inst/LUT__4934  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .I3(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n3340 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fb8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4934 .LUTMASK = 16'h0fb8;
    EFX_LUT4 \edb_top_inst/LUT__4935  (.I0(\edb_top_inst/n3340 ), .I1(jtag_inst2_SEL), 
            .I2(jtag_inst2_UPDATE), .I3(\edb_top_inst/edb_user_dr[81] ), 
            .O(\edb_top_inst/debug_hub_inst/n266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4935 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4936  (.I0(jtag_inst2_SEL), .I1(jtag_inst2_SHIFT), 
            .O(\edb_top_inst/debug_hub_inst/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4936 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4937  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[3] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[1] ), .O(\edb_top_inst/n2739 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4937 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4945  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4945 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4946  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4946 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4947  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4947 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4948  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4948 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4949  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4949 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4950  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4950 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4951  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4951 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4952  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4952 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4953  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4953 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4954  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4954 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4955  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4955 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4956  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4956 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4957  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4957 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4958  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4958 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4959  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4959 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4960  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4960 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4961  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4961 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4962  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4962 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4963  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4963 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4964  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4964 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4965  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4965 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4966  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4966 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4967  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4967 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4968  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4968 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4969  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4969 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4970  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4970 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4971  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4971 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4972  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4972 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4973  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i35_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4973 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4974  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i36_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4974 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4975  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i37_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4975 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4976  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i38_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4976 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4977  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i39_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4977 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4978  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i40_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4978 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__3984  (.I0(\edb_top_inst/la0/crc_data_out[21] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/la0/crc_data_out[22] ), 
            .I3(\edb_top_inst/edb_user_dr[72] ), .O(\edb_top_inst/n2758 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3984 .LUTMASK = 16'h9009;
    EFX_ADD \edb_top_inst/la0/add_91/i1  (.I0(\edb_top_inst/la0/address_counter[0] ), 
            .I1(\edb_top_inst/n1249 ), .CI(1'b0), .O(\edb_top_inst/n67 ), 
            .CO(\edb_top_inst/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i2  (.I0(\edb_top_inst/la0/bit_count[1] ), 
            .I1(\edb_top_inst/la0/bit_count[0] ), .CI(1'b0), .O(\edb_top_inst/n69 ), 
            .CO(\edb_top_inst/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_100/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .CI(1'b0), 
            .O(\edb_top_inst/n73 ), .CO(\edb_top_inst/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
            .CI(1'b0), .O(\edb_top_inst/n693 ), .CO(\edb_top_inst/n694 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
            .CI(1'b0), .O(\edb_top_inst/n695 ), .CO(\edb_top_inst/n696 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .CI(1'b0), 
            .CO(\edb_top_inst/n697 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_sample_cnt[0] ), .CI(1'b0), .CO(\edb_top_inst/n698 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(1'b1), .CI(n10138), .O(\edb_top_inst/n710 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4673)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I1(1'b1), .CI(n10139), .O(\edb_top_inst/n711 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4659)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i13  (.I0(\edb_top_inst/la0/la_sample_cnt[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n714 ), .O(\edb_top_inst/n712 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12  (.I0(\edb_top_inst/la0/la_sample_cnt[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n716 ), .O(\edb_top_inst/n713 ), 
            .CO(\edb_top_inst/n714 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11  (.I0(\edb_top_inst/la0/la_sample_cnt[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n718 ), .O(\edb_top_inst/n715 ), 
            .CO(\edb_top_inst/n716 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10  (.I0(\edb_top_inst/la0/la_sample_cnt[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n720 ), .O(\edb_top_inst/n717 ), 
            .CO(\edb_top_inst/n718 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9  (.I0(\edb_top_inst/la0/la_sample_cnt[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n722 ), .O(\edb_top_inst/n719 ), 
            .CO(\edb_top_inst/n720 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8  (.I0(\edb_top_inst/la0/la_sample_cnt[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n724 ), .O(\edb_top_inst/n721 ), 
            .CO(\edb_top_inst/n722 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7  (.I0(\edb_top_inst/la0/la_sample_cnt[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n726 ), .O(\edb_top_inst/n723 ), 
            .CO(\edb_top_inst/n724 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6  (.I0(\edb_top_inst/la0/la_sample_cnt[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n728 ), .O(\edb_top_inst/n725 ), 
            .CO(\edb_top_inst/n726 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5  (.I0(\edb_top_inst/la0/la_sample_cnt[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n730 ), .O(\edb_top_inst/n727 ), 
            .CO(\edb_top_inst/n728 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4  (.I0(\edb_top_inst/la0/la_sample_cnt[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n732 ), .O(\edb_top_inst/n729 ), 
            .CO(\edb_top_inst/n730 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3  (.I0(\edb_top_inst/la0/la_sample_cnt[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n698 ), .O(\edb_top_inst/n731 ), 
            .CO(\edb_top_inst/n732 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i13  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n735 ), .O(\edb_top_inst/n733 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n737 ), .O(\edb_top_inst/n734 ), 
            .CO(\edb_top_inst/n735 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n739 ), .O(\edb_top_inst/n736 ), 
            .CO(\edb_top_inst/n737 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n741 ), .O(\edb_top_inst/n738 ), 
            .CO(\edb_top_inst/n739 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n743 ), .O(\edb_top_inst/n740 ), 
            .CO(\edb_top_inst/n741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n745 ), .O(\edb_top_inst/n742 ), 
            .CO(\edb_top_inst/n743 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n747 ), .O(\edb_top_inst/n744 ), 
            .CO(\edb_top_inst/n745 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n749 ), .O(\edb_top_inst/n746 ), 
            .CO(\edb_top_inst/n747 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n751 ), .O(\edb_top_inst/n748 ), 
            .CO(\edb_top_inst/n749 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n753 ), .O(\edb_top_inst/n750 ), 
            .CO(\edb_top_inst/n751 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n697 ), .O(\edb_top_inst/n752 ), 
            .CO(\edb_top_inst/n753 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i12  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n841 ), .O(\edb_top_inst/n838 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n843 ), .O(\edb_top_inst/n840 ), 
            .CO(\edb_top_inst/n841 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n845 ), .O(\edb_top_inst/n842 ), 
            .CO(\edb_top_inst/n843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n847 ), .O(\edb_top_inst/n844 ), 
            .CO(\edb_top_inst/n845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n849 ), .O(\edb_top_inst/n846 ), 
            .CO(\edb_top_inst/n847 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n851 ), .O(\edb_top_inst/n848 ), 
            .CO(\edb_top_inst/n849 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n853 ), .O(\edb_top_inst/n850 ), 
            .CO(\edb_top_inst/n851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n855 ), .O(\edb_top_inst/n852 ), 
            .CO(\edb_top_inst/n853 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n857 ), .O(\edb_top_inst/n854 ), 
            .CO(\edb_top_inst/n855 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n696 ), .O(\edb_top_inst/n856 ), 
            .CO(\edb_top_inst/n857 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i12  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1009 ), .O(\edb_top_inst/n1005 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1012 ), .O(\edb_top_inst/n1008 ), 
            .CO(\edb_top_inst/n1009 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1014 ), .O(\edb_top_inst/n1011 ), 
            .CO(\edb_top_inst/n1012 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1016 ), .O(\edb_top_inst/n1013 ), 
            .CO(\edb_top_inst/n1014 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1018 ), .O(\edb_top_inst/n1015 ), 
            .CO(\edb_top_inst/n1016 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1020 ), .O(\edb_top_inst/n1017 ), 
            .CO(\edb_top_inst/n1018 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1022 ), .O(\edb_top_inst/n1019 ), 
            .CO(\edb_top_inst/n1020 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1024 ), .O(\edb_top_inst/n1021 ), 
            .CO(\edb_top_inst/n1022 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1026 ), .O(\edb_top_inst/n1023 ), 
            .CO(\edb_top_inst/n1024 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n694 ), .O(\edb_top_inst/n1025 ), 
            .CO(\edb_top_inst/n1026 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i12  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1029 ), .O(\edb_top_inst/n1027 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1031 ), .O(\edb_top_inst/n1028 ), 
            .CO(\edb_top_inst/n1029 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1033 ), .O(\edb_top_inst/n1030 ), 
            .CO(\edb_top_inst/n1031 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1035 ), .O(\edb_top_inst/n1032 ), 
            .CO(\edb_top_inst/n1033 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1037 ), .O(\edb_top_inst/n1034 ), 
            .CO(\edb_top_inst/n1035 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1039 ), .O(\edb_top_inst/n1036 ), 
            .CO(\edb_top_inst/n1037 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1041 ), .O(\edb_top_inst/n1038 ), 
            .CO(\edb_top_inst/n1039 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1043 ), .O(\edb_top_inst/n1040 ), 
            .CO(\edb_top_inst/n1041 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1045 ), .O(\edb_top_inst/n1042 ), 
            .CO(\edb_top_inst/n1043 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n74 ), .O(\edb_top_inst/n1044 ), 
            .CO(\edb_top_inst/n1045 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i6  (.I0(\edb_top_inst/la0/bit_count[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1048 ), .O(\edb_top_inst/n1046 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_100/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i5  (.I0(\edb_top_inst/la0/bit_count[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1050 ), .O(\edb_top_inst/n1047 ), 
            .CO(\edb_top_inst/n1048 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_100/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i4  (.I0(\edb_top_inst/la0/bit_count[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1052 ), .O(\edb_top_inst/n1049 ), 
            .CO(\edb_top_inst/n1050 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_100/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i3  (.I0(\edb_top_inst/la0/bit_count[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n70 ), .O(\edb_top_inst/n1051 ), 
            .CO(\edb_top_inst/n1052 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_100/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i27  (.I0(\edb_top_inst/la0/address_counter[26] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1065 ), .O(\edb_top_inst/n1062 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i27 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i26  (.I0(\edb_top_inst/la0/address_counter[25] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1067 ), .O(\edb_top_inst/n1064 ), 
            .CO(\edb_top_inst/n1065 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i26 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i25  (.I0(\edb_top_inst/la0/address_counter[24] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1069 ), .O(\edb_top_inst/n1066 ), 
            .CO(\edb_top_inst/n1067 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i25 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i24  (.I0(\edb_top_inst/la0/address_counter[23] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1071 ), .O(\edb_top_inst/n1068 ), 
            .CO(\edb_top_inst/n1069 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i24 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i23  (.I0(\edb_top_inst/la0/address_counter[22] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1073 ), .O(\edb_top_inst/n1070 ), 
            .CO(\edb_top_inst/n1071 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i23 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i22  (.I0(\edb_top_inst/la0/address_counter[21] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1075 ), .O(\edb_top_inst/n1072 ), 
            .CO(\edb_top_inst/n1073 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i22 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i21  (.I0(\edb_top_inst/la0/address_counter[20] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1077 ), .O(\edb_top_inst/n1074 ), 
            .CO(\edb_top_inst/n1075 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i21 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i20  (.I0(\edb_top_inst/la0/address_counter[19] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1079 ), .O(\edb_top_inst/n1076 ), 
            .CO(\edb_top_inst/n1077 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i20 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i19  (.I0(\edb_top_inst/la0/address_counter[18] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1081 ), .O(\edb_top_inst/n1078 ), 
            .CO(\edb_top_inst/n1079 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i19 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i18  (.I0(\edb_top_inst/la0/address_counter[17] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1083 ), .O(\edb_top_inst/n1080 ), 
            .CO(\edb_top_inst/n1081 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i18 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i17  (.I0(\edb_top_inst/la0/address_counter[16] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1085 ), .O(\edb_top_inst/n1082 ), 
            .CO(\edb_top_inst/n1083 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i17 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i16  (.I0(\edb_top_inst/la0/address_counter[15] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1087 ), .O(\edb_top_inst/n1084 ), 
            .CO(\edb_top_inst/n1085 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i16 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i15  (.I0(\edb_top_inst/la0/address_counter[14] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1089 ), .O(\edb_top_inst/n1086 ), 
            .CO(\edb_top_inst/n1087 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i15 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i14  (.I0(\edb_top_inst/la0/address_counter[13] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1091 ), .O(\edb_top_inst/n1088 ), 
            .CO(\edb_top_inst/n1089 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i13  (.I0(\edb_top_inst/la0/address_counter[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1093 ), .O(\edb_top_inst/n1090 ), 
            .CO(\edb_top_inst/n1091 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i12  (.I0(\edb_top_inst/la0/address_counter[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1095 ), .O(\edb_top_inst/n1092 ), 
            .CO(\edb_top_inst/n1093 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i11  (.I0(\edb_top_inst/la0/address_counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1097 ), .O(\edb_top_inst/n1094 ), 
            .CO(\edb_top_inst/n1095 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i10  (.I0(\edb_top_inst/la0/address_counter[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1099 ), .O(\edb_top_inst/n1096 ), 
            .CO(\edb_top_inst/n1097 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i9  (.I0(\edb_top_inst/la0/address_counter[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1101 ), .O(\edb_top_inst/n1098 ), 
            .CO(\edb_top_inst/n1099 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i8  (.I0(\edb_top_inst/la0/address_counter[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1103 ), .O(\edb_top_inst/n1100 ), 
            .CO(\edb_top_inst/n1101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i7  (.I0(\edb_top_inst/la0/address_counter[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1105 ), .O(\edb_top_inst/n1102 ), 
            .CO(\edb_top_inst/n1103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i6  (.I0(\edb_top_inst/la0/address_counter[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1107 ), .O(\edb_top_inst/n1104 ), 
            .CO(\edb_top_inst/n1105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i5  (.I0(\edb_top_inst/la0/address_counter[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1109 ), .O(\edb_top_inst/n1106 ), 
            .CO(\edb_top_inst/n1107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i4  (.I0(\edb_top_inst/la0/address_counter[3] ), 
            .I1(\edb_top_inst/n2733 ), .CI(\edb_top_inst/n1111 ), .O(\edb_top_inst/n1108 ), 
            .CO(\edb_top_inst/n1109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i3  (.I0(\edb_top_inst/la0/address_counter[2] ), 
            .I1(\edb_top_inst/n2736 ), .CI(\edb_top_inst/n1113 ), .O(\edb_top_inst/n1110 ), 
            .CO(\edb_top_inst/n1111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i2  (.I0(\edb_top_inst/la0/address_counter[1] ), 
            .I1(\edb_top_inst/n2739 ), .CI(\edb_top_inst/n68 ), .O(\edb_top_inst/n1112 ), 
            .CO(\edb_top_inst/n1113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i12  (.I0(\edb_top_inst/la0/address_counter[26] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1126 ), .O(\edb_top_inst/n1123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i11  (.I0(\edb_top_inst/la0/address_counter[25] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1128 ), .O(\edb_top_inst/n1125 ), 
            .CO(\edb_top_inst/n1126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i10  (.I0(\edb_top_inst/la0/address_counter[24] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1130 ), .O(\edb_top_inst/n1127 ), 
            .CO(\edb_top_inst/n1128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i9  (.I0(\edb_top_inst/la0/address_counter[23] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1132 ), .O(\edb_top_inst/n1129 ), 
            .CO(\edb_top_inst/n1130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i8  (.I0(\edb_top_inst/la0/address_counter[22] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1134 ), .O(\edb_top_inst/n1131 ), 
            .CO(\edb_top_inst/n1132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i7  (.I0(\edb_top_inst/la0/address_counter[21] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1136 ), .O(\edb_top_inst/n1133 ), 
            .CO(\edb_top_inst/n1134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i6  (.I0(\edb_top_inst/la0/address_counter[20] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1138 ), .O(\edb_top_inst/n1135 ), 
            .CO(\edb_top_inst/n1136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i5  (.I0(\edb_top_inst/la0/address_counter[19] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1143 ), .O(\edb_top_inst/n1137 ), 
            .CO(\edb_top_inst/n1138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i4  (.I0(\edb_top_inst/la0/address_counter[18] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1145 ), .O(\edb_top_inst/n1142 ), 
            .CO(\edb_top_inst/n1143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i3  (.I0(\edb_top_inst/la0/address_counter[17] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1147 ), .O(\edb_top_inst/n1144 ), 
            .CO(\edb_top_inst/n1145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i2  (.I0(\edb_top_inst/la0/address_counter[16] ), 
            .I1(\edb_top_inst/la0/address_counter[15] ), .CI(1'b0), .O(\edb_top_inst/n1146 ), 
            .CO(\edb_top_inst/n1147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i2 .I1_POLARITY = 1'b1;
    EFX_LUT4 LUT__13630 (.I0(\MCsiRxController/MCsi2Decoder/wFtiRd[16] ), 
            .I1(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), .I2(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), 
            .I3(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .O(\MCsiRxController/MCsi2Decoder/n630 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h03e0 */ ;
    defparam LUT__13630.LUTMASK = 16'h03e0;
    EFX_LUT4 LUT__13631 (.I0(rSRST), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), 
            .O(\MCsiRxController/MCsi2Decoder/n632 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__13631.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__13632 (.I0(oTestPort[24]), .I1(oTestPort[0]), .O(\MCsiRxController/MCsi2Decoder/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__13632.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__13633 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
            .O(n9759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13633.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13634 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] ), 
            .O(n9760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13634.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13635 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
            .O(n9761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13635.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13636 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] ), 
            .O(n9762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13636.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13637 (.I0(n9759), .I1(n9760), .I2(n9761), .I3(n9762), 
            .O(n9763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13637.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13638 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
            .O(n9764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13638.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13639 (.I0(n9763), .I1(n9764), .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRVd )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777 */ ;
    defparam LUT__13639.LUTMASK = 16'h7777;
    EFX_LUT4 LUT__13640 (.I0(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), .O(n9765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__13640.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__13641 (.I0(\wHsDatatype[2] ), .I1(\wHsDatatype[3] ), .I2(\wHsDatatype[4] ), 
            .I3(\wHsDatatype[5] ), .O(n9766)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__13641.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__13642 (.I0(n9766), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .I3(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), 
            .O(n9767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__13642.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__13643 (.I0(n9767), .I1(n9765), .I2(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), 
            .O(\~MCsiRxController/MCsi2Decoder/reduce_nor_75/n1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f1f */ ;
    defparam LUT__13643.LUTMASK = 16'h1f1f;
    EFX_LUT4 LUT__13644 (.I0(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), .I3(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), 
            .O(\MCsiRxController/MCsi2Decoder/n603 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1800 */ ;
    defparam LUT__13644.LUTMASK = 16'h1800;
    EFX_LUT4 LUT__13645 (.I0(\wHsWordCnt[1] ), .I1(\wHsWordCnt[2] ), .I2(\wHsWordCnt[3] ), 
            .I3(\wHsWordCnt[4] ), .O(n9768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13645.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13646 (.I0(\wHsWordCnt[6] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5] ), 
            .O(n9769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__13646.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__13647 (.I0(\wHsWordCnt[5] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4] ), 
            .I2(n9768), .I3(n9769), .O(n9770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd6bf */ ;
    defparam LUT__13647.LUTMASK = 16'hd6bf;
    EFX_LUT4 LUT__13648 (.I0(\wHsWordCnt[5] ), .I1(\wHsWordCnt[6] ), .I2(\wHsWordCnt[7] ), 
            .I3(\wHsWordCnt[8] ), .O(n9771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13648.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13649 (.I0(\wHsWordCnt[9] ), .I1(n9768), .I2(n9771), 
            .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9] ), .O(n9772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40bf */ ;
    defparam LUT__13649.LUTMASK = 16'h40bf;
    EFX_LUT4 LUT__13650 (.I0(\wHsWordCnt[7] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6] ), 
            .I2(\wHsWordCnt[8] ), .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7] ), 
            .O(n9773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13650.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13651 (.I0(\wHsWordCnt[7] ), .I1(\wHsWordCnt[8] ), .I2(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7] ), 
            .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6] ), .O(n9774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d */ ;
    defparam LUT__13651.LUTMASK = 16'heb7d;
    EFX_LUT4 LUT__13652 (.I0(n9774), .I1(n9773), .I2(\wHsWordCnt[6] ), 
            .I3(n9769), .O(n9775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h333a */ ;
    defparam LUT__13652.LUTMASK = 16'h333a;
    EFX_LUT4 LUT__13653 (.I0(\wHsWordCnt[11] ), .I1(\wHsWordCnt[12] ), .I2(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] ), 
            .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] ), .O(n9776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d */ ;
    defparam LUT__13653.LUTMASK = 16'heb7d;
    EFX_LUT4 LUT__13654 (.I0(\wHsWordCnt[11] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] ), 
            .I2(\wHsWordCnt[12] ), .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] ), 
            .O(n9777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13654.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13655 (.I0(n9776), .I1(n9777), .I2(\wHsWordCnt[10] ), 
            .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9] ), .O(n9778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a33 */ ;
    defparam LUT__13655.LUTMASK = 16'h3a33;
    EFX_LUT4 LUT__13656 (.I0(n9775), .I1(n9778), .I2(n9772), .I3(\wHsWordCnt[10] ), 
            .O(n9779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110 */ ;
    defparam LUT__13656.LUTMASK = 16'h0110;
    EFX_LUT4 LUT__13657 (.I0(\wHsWordCnt[9] ), .I1(\wHsWordCnt[10] ), .I2(\wHsWordCnt[11] ), 
            .I3(\wHsWordCnt[12] ), .O(n9780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13657.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13658 (.I0(n9768), .I1(n9771), .I2(n9780), .O(n9781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13658.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13659 (.I0(\wHsWordCnt[14] ), .I1(n9781), .I2(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12] ), 
            .I3(\wHsWordCnt[13] ), .O(n9782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7e */ ;
    defparam LUT__13659.LUTMASK = 16'heb7e;
    EFX_LUT4 LUT__13660 (.I0(\wHsWordCnt[4] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3] ), 
            .O(n9783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__13660.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__13661 (.I0(\wHsWordCnt[1] ), .I1(\wHsWordCnt[2] ), .O(n9784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13661.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13662 (.I0(\wHsWordCnt[3] ), .I1(n9783), .I2(n9784), 
            .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2] ), .O(n9785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__13662.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__13663 (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] ), 
            .I1(\wHsWordCnt[2] ), .I2(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1] ), 
            .I3(\wHsWordCnt[1] ), .O(n9786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbed7 */ ;
    defparam LUT__13663.LUTMASK = 16'hbed7;
    EFX_LUT4 LUT__13664 (.I0(n9786), .I1(\wHsWordCnt[15] ), .I2(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), 
            .O(n9787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__13664.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__13665 (.I0(n9768), .I1(n9771), .I2(\wHsWordCnt[9] ), 
            .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8] ), .O(n9788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7887 */ ;
    defparam LUT__13665.LUTMASK = 16'h7887;
    EFX_LUT4 LUT__13666 (.I0(n9785), .I1(n9787), .I2(n9788), .O(n9789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__13666.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__13667 (.I0(n9770), .I1(n9782), .I2(n9779), .I3(n9789), 
            .O(n9790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__13667.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__13668 (.I0(n9790), .I1(rSRST), .O(\MCsiRxController/MCsi2Decoder/qLineCntRst )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__13668.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__13669 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .O(n9791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13669.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13670 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .O(n9792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13670.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13671 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .O(n9793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13671.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13672 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .O(n9794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13672.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13673 (.I0(n9791), .I1(n9792), .I2(n9793), .I3(n9794), 
            .O(n9795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13673.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13674 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] ), 
            .O(n9796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13674.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13675 (.I0(n9795), .I1(n9796), .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/equal_38/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777 */ ;
    defparam LUT__13675.LUTMASK = 16'h7777;
    EFX_LUT4 LUT__13676 (.I0(\MCsiRxController/MCsi2Decoder/wFtiEmp[0] ), 
            .I1(wCdcFifoFull), .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/equal_38/n19 ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__13676.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__13677 (.I0(n9790), .I1(n9765), .I2(n9767), .O(\MCsiRxController/MCsi2Decoder/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__13677.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__13678 (.I0(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), .I2(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), 
            .O(\MCsiRxController/MCsi2Decoder/n606 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2c2c */ ;
    defparam LUT__13678.LUTMASK = 16'h2c2c;
    EFX_LUT4 LUT__13679 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n233 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13679.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13680 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n238 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13680.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13681 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n243 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__13681.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__13682 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .O(n9797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13682.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13683 (.I0(n9797), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13683.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13684 (.I0(n9797), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n253 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13684.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13685 (.I0(n9797), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n258 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__13685.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__13686 (.I0(n9797), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] ), 
            .O(n9798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13686.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13687 (.I0(n9798), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n263 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13687.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13688 (.I0(n9798), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n268 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13688.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13689 (.I0(n9798), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n273 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__13689.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__13690 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .O(n9799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13690.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13691 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] ), 
            .O(n9800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13691.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13692 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .O(n9801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13692.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13693 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .O(n9802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13693.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13694 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .O(n9803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13694.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13695 (.I0(n9800), .I1(n9801), .I2(n9802), .I3(n9803), 
            .O(n9804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13695.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13696 (.I0(n9804), .I1(n9799), .I2(\MCsiRxController/MCsi2Decoder/wFtiEmp[0] ), 
            .I3(wCdcFifoFull), .O(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__13696.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__13697 (.I0(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .O(\MCsiRxController/MCsi2Decoder/equal_62/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__13697.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__13698 (.I0(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), .O(\MCsiRxController/MCsi2Decoder/equal_59/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__13698.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__13699 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] ), .O(n9805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__13699.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__13700 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] ), .O(n9806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__13700.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__13701 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] ), .O(n9807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13701.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13702 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), .O(n9808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13702.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13703 (.I0(n9808), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), .O(n9809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141 */ ;
    defparam LUT__13703.LUTMASK = 16'h4141;
    EFX_LUT4 LUT__13704 (.I0(n9807), .I1(n9806), .I2(n9805), .I3(n9809), 
            .O(n9810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__13704.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__13705 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .O(n9811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13705.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13706 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .O(n9812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13706.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13707 (.I0(n9810), .I1(n9811), .I2(n9812), .O(\MCsiRxController/genblk1[0].mVideoFIFO/equal_75/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f7f */ ;
    defparam LUT__13707.LUTMASK = 16'h7f7f;
    EFX_LUT4 LUT__13708 (.I0(\MCsiRxController/wFtiEmp[0] ), .I1(wVideofull), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/equal_75/n17 ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__13708.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__13709 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), .O(n9813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__13709.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__13710 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), .O(n9814)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13710.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13711 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .I2(n9814), 
            .O(n9815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__13711.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__13712 (.I0(n9811), .I1(n9813), .I2(n9815), .O(n9816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__13712.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__13713 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] ), .O(n9817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13713.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13714 (.I0(n9817), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] ), .O(n9818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13714.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13715 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
            .I1(n9806), .I2(n9818), .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] ), 
            .O(n9819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__13715.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__13716 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), .I2(n9805), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .O(n9820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f */ ;
    defparam LUT__13716.LUTMASK = 16'hed3f;
    EFX_LUT4 LUT__13717 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] ), .O(n9821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13717.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13718 (.I0(n9817), .I1(n9821), .I2(n9808), .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), 
            .O(n9822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6ffc */ ;
    defparam LUT__13718.LUTMASK = 16'h6ffc;
    EFX_LUT4 LUT__13719 (.I0(n9819), .I1(n9820), .I2(n9822), .O(n9823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__13719.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__13720 (.I0(n9805), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), .O(n9824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7e7 */ ;
    defparam LUT__13720.LUTMASK = 16'he7e7;
    EFX_LUT4 LUT__13721 (.I0(n9824), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), .O(n9825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141 */ ;
    defparam LUT__13721.LUTMASK = 16'h4141;
    EFX_LUT4 LUT__13722 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
            .I1(n9807), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] ), 
            .I3(n9806), .O(n9826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc8bf */ ;
    defparam LUT__13722.LUTMASK = 16'hc8bf;
    EFX_LUT4 LUT__13723 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
            .I1(n9807), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] ), 
            .I3(n9817), .O(n9827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde */ ;
    defparam LUT__13723.LUTMASK = 16'hbdde;
    EFX_LUT4 LUT__13724 (.I0(n9826), .I1(n9827), .I2(n9825), .I3(n9816), 
            .O(n9828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__13724.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__13725 (.I0(n9810), .I1(n9816), .I2(n9823), .I3(n9828), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/qFullAllmost )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff2 */ ;
    defparam LUT__13725.LUTMASK = 16'hfff2;
    EFX_LUT4 LUT__13726 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[4] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[7] ), .O(n9829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13726.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13727 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[0] ), .I2(n9829), 
            .O(n9830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__13727.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__13728 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[2] ), .O(n9831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13728.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13729 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[3] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[6] ), .O(n9832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13729.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13730 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[5] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[8] ), .O(n9833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13730.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13731 (.I0(n9830), .I1(n9831), .I2(n9832), .I3(n9833), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/qRVD )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__13731.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__13732 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/n436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13732.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13733 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/n441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13733.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13734 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/n446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__13734.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__13735 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .O(n9834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13735.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13736 (.I0(n9834), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/n451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13736.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13737 (.I0(n9834), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/n456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13737.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13738 (.I0(n9817), .I1(n9834), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] ), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/n461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13738.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13739 (.I0(n9817), .I1(n9834), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/n466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__13739.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__13740 (.I0(n9817), .I1(n9834), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] ), .O(n9835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13740.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13741 (.I0(n9835), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] ), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/n471 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13741.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13742 (.I0(oTestPort[24]), .I1(n3828), .O(\MCsiRxController/n278 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13742.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13743 (.I0(oTestPort[24]), .I1(n3826), .O(\MCsiRxController/n277 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13743.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13744 (.I0(oTestPort[24]), .I1(n3824), .O(\MCsiRxController/n276 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13744.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13745 (.I0(oTestPort[24]), .I1(n3822), .O(\MCsiRxController/n275 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13745.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13746 (.I0(oTestPort[24]), .I1(n3820), .O(\MCsiRxController/n274 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13746.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13747 (.I0(oTestPort[24]), .I1(n3818), .O(\MCsiRxController/n273 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13747.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13748 (.I0(oTestPort[24]), .I1(n3816), .O(\MCsiRxController/n272 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13748.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13749 (.I0(oTestPort[24]), .I1(n3814), .O(\MCsiRxController/n271 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13749.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13750 (.I0(oTestPort[24]), .I1(n3812), .O(\MCsiRxController/n270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13750.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13751 (.I0(oTestPort[24]), .I1(n3810), .O(\MCsiRxController/n269 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13751.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13752 (.I0(oTestPort[24]), .I1(n3808), .O(\MCsiRxController/n268 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13752.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13753 (.I0(oTestPort[24]), .I1(n3806), .O(\MCsiRxController/n267 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13753.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13754 (.I0(oTestPort[24]), .I1(n3804), .O(\MCsiRxController/n266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13754.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13755 (.I0(oTestPort[24]), .I1(n3802), .O(\MCsiRxController/n265 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13755.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13756 (.I0(oTestPort[24]), .I1(n3801), .O(\MCsiRxController/n264 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13756.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13757 (.I0(wVideoVd), .I1(\MVideoPostProcess/rVtgRstSel ), 
            .O(\MVideoPostProcess/qVtgRstCntCke )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13757.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13758 (.I0(\MVideoPostProcess/rVtgRstCnt[8] ), .I1(\MVideoPostProcess/rVtgRstCnt[9] ), 
            .I2(\MVideoPostProcess/rVtgRstCnt[10] ), .O(n9836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13758.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13759 (.I0(\MVideoPostProcess/rVtgRstCnt[4] ), .I1(\MVideoPostProcess/rVtgRstCnt[5] ), 
            .I2(\MVideoPostProcess/rVtgRstCnt[6] ), .I3(\MVideoPostProcess/rVtgRstCnt[7] ), 
            .O(n9837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__13759.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__13760 (.I0(\MVideoPostProcess/rVtgRstCnt[0] ), .I1(\MVideoPostProcess/rVtgRstCnt[1] ), 
            .I2(\MVideoPostProcess/rVtgRstCnt[2] ), .I3(\MVideoPostProcess/rVtgRstCnt[3] ), 
            .O(n9838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13760.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13761 (.I0(n9836), .I1(n9837), .I2(n9838), .O(\MVideoPostProcess/equal_18/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f7f */ ;
    defparam LUT__13761.LUTMASK = 16'h7f7f;
    EFX_LUT4 LUT__13762 (.I0(\MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\~n1834 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13762.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13763 (.I0(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0] ), 
            .O(n9839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__13763.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__13764 (.I0(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] ), 
            .I3(n9839), .O(n9840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__13764.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__13765 (.I0(n9840), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] ), .O(n9841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13765.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13766 (.I0(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_ack ), .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(n9842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__13766.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__13767 (.I0(n9841), .I1(n9842), .O(n9843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13767.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13768 (.I0(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .I1(pll_inst1_LOCKED), .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I3(rBRST), .O(n9844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__13768.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__13769 (.I0(n9843), .I1(n9844), .O(ceg_net939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__13769.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__13770 (.I0(\MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] ), 
            .I1(n9841), .I2(n9842), .O(\MVideoPostProcess/inst_adv7511_config/n816 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f1f */ ;
    defparam LUT__13770.LUTMASK = 16'h1f1f;
    EFX_LUT4 LUT__13771 (.I0(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3] ), .O(n9845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13771.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13772 (.I0(n9845), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6] ), 
            .O(n9846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13772.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13773 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_2P ), 
            .I1(n9846), .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_3P ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7] ), .O(n9847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__13773.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__13774 (.I0(n9847), .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .I3(n9844), .O(\~ceg_net512 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__13774.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__13775 (.I0(n9843), .I1(\MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n833 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13775.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13776 (.I0(\MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n268 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13776.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13777 (.I0(\MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] ), 
            .I1(n9843), .I2(n9844), .O(ceg_net995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f8f */ ;
    defparam LUT__13777.LUTMASK = 16'h8f8f;
    EFX_LUT4 LUT__13778 (.I0(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n1107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13778.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13779 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_2P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/n1107 ), .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_3P ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n1224 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__13779.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__13780 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n277 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__13780.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__13781 (.I0(rBRST), .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(ceg_net479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__13781.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__13782 (.I0(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n242 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13782.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13783 (.I0(ceg_net479), .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(n9848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13783.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13784 (.I0(\MVideoPostProcess/inst_adv7511_config/w_ack ), 
            .I1(n9841), .I2(n9848), .I3(\~ceg_net512 ), .O(ceg_net1327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__13784.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__13785 (.I0(rBRST), .I1(\MVideoPostProcess/inst_adv7511_config/n1107 ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n1243 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13785.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13786 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .O(n9849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13786.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13787 (.I0(iAdv7511Scl), .I1(oAdv7511SclOe), .I2(n9849), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), .O(n9850)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__13787.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__13788 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n9851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13788.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13789 (.I0(n9850), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I3(n9851), .O(n9852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe0f */ ;
    defparam LUT__13789.LUTMASK = 16'hfe0f;
    EFX_LUT4 LUT__13790 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(n9852), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n846 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13790.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13791 (.I0(n9851), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n9853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13791.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13792 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] ), 
            .I1(n9853), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n852 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13792.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13793 (.I0(n9849), .I1(iAdv7511Sda), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n9854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__13793.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__13794 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I1(n9849), .O(n9855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13794.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13795 (.I0(n9854), .I1(n9855), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I3(n9851), .O(ceg_net1087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe03 */ ;
    defparam LUT__13795.LUTMASK = 16'hfe03;
    EFX_LUT4 LUT__13796 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n9856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13796.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13797 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2] ), 
            .O(n9857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13797.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13798 (.I0(\MVideoPostProcess/inst_adv7511_config/r_last_1P ), 
            .I1(oAdv7511SdaOe), .I2(n9849), .I3(n9857), .O(n9858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccc */ ;
    defparam LUT__13798.LUTMASK = 16'h5ccc;
    EFX_LUT4 LUT__13799 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), .I2(oAdv7511SdaOe), 
            .I3(n9849), .O(n9859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__13799.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__13800 (.I0(n9859), .I1(n9858), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n9860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__13800.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__13801 (.I0(iAdv7511Sda), .I1(oAdv7511SdaOe), .O(n9861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__13801.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__13802 (.I0(n9857), .I1(n9861), .O(n9862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13802.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13803 (.I0(n9862), .I1(n9849), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] ), 
            .O(n9863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__13803.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__13804 (.I0(iAdv7511Sda), .I1(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
            .O(n9864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13804.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13805 (.I0(n9849), .I1(oAdv7511SdaOe), .I2(n9864), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n9865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__13805.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__13806 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(n9856), .O(n9866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13806.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13807 (.I0(iAdv7511Sda), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(n9866), .O(n9867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__13807.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__13808 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n9868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13808.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13809 (.I0(n9868), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n9869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13809.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13810 (.I0(n9867), .I1(n9869), .I2(n9863), .I3(n9865), 
            .O(n9870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__13810.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__13811 (.I0(n9849), .I1(n9851), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n9871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__13811.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__13812 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(n9851), .O(n9872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13812.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13813 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] ), 
            .I1(iAdv7511Sda), .I2(n9849), .I3(n9872), .O(n9873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__13813.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__13814 (.I0(n9873), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(oAdv7511SdaOe), .I3(n9871), .O(n9874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__13814.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__13815 (.I0(n9860), .I1(n9856), .I2(n9870), .I3(n9874), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n847 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8ff */ ;
    defparam LUT__13815.LUTMASK = 16'hf8ff;
    EFX_LUT4 LUT__13816 (.I0(iAdv7511Scl), .I1(oAdv7511SclOe), .I2(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
            .I3(n9849), .O(n9875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__13816.LUTMASK = 16'he000;
    EFX_LUT4 LUT__13817 (.I0(n9849), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n9876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13817.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13818 (.I0(n9875), .I1(n9876), .I2(n9872), .O(ceg_net566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__13818.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__13819 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(ceg_net566), .O(n9877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__13819.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__13820 (.I0(n9849), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n9878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__13820.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__13821 (.I0(n9849), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(n9866), .I3(n9878), .O(n9879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__13821.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__13822 (.I0(n9877), .I1(n9879), .O(ceg_net1335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__13822.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__13823 (.I0(iAdv7511Sda), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n9880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfcc4 */ ;
    defparam LUT__13823.LUTMASK = 16'hfcc4;
    EFX_LUT4 LUT__13824 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .I1(n9861), .I2(n9851), .I3(n9880), .O(n9881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__13824.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__13825 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(n9881), .I2(n9871), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n848 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f1 */ ;
    defparam LUT__13825.LUTMASK = 16'h00f1;
    EFX_LUT4 LUT__13826 (.I0(n9849), .I1(n9857), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n9882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13826.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13827 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I1(n9875), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I3(n9851), .O(n9883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb0f */ ;
    defparam LUT__13827.LUTMASK = 16'hfb0f;
    EFX_LUT4 LUT__13828 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I1(n9882), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .I3(n9883), .O(ceg_net1400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__13828.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__13829 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n870 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13829.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13830 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I1(n9861), .I2(n9857), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n9884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__13830.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__13831 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .I1(n9864), .I2(n9849), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n9885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__13831.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__13832 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n9886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbaa3 */ ;
    defparam LUT__13832.LUTMASK = 16'hbaa3;
    EFX_LUT4 LUT__13833 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0] ), 
            .I1(n9885), .I2(n9866), .I3(n9886), .O(n9887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__13833.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__13834 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0] ), 
            .I1(n9884), .I2(n9868), .I3(n9887), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n879 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__13834.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__13835 (.I0(n9864), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n9888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13835.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13836 (.I0(n9849), .I1(n9866), .I2(n9872), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n9889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__13836.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__13837 (.I0(n9888), .I1(n9849), .I2(n9869), .I3(n9889), 
            .O(ceg_net1463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffb0 */ ;
    defparam LUT__13837.LUTMASK = 16'hffb0;
    EFX_LUT4 LUT__13842 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n9892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13842.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13843 (.I0(n9864), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n9893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13843.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13844 (.I0(n9892), .I1(iAdv7511Sda), .I2(n9893), .I3(n9868), 
            .O(n9894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__13844.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__13845 (.I0(n9862), .I1(n9849), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n9895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__13845.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__13846 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(n9861), .O(n9896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13846.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13847 (.I0(n9896), .I1(n9857), .I2(n9856), .O(n9897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__13847.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__13848 (.I0(n9897), .I1(n9851), .I2(n9855), .O(n9898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__13848.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__13849 (.I0(n9849), .I1(iAdv7511Sda), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n9899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;
    defparam LUT__13849.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__13850 (.I0(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .I2(n9899), .O(n9900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__13850.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__13851 (.I0(n9900), .I1(n9856), .I2(n9871), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n9901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__13851.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__13852 (.I0(n9895), .I1(n9894), .I2(n9898), .I3(n9901), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n829 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4 */ ;
    defparam LUT__13852.LUTMASK = 16'hfff4;
    EFX_LUT4 LUT__13853 (.I0(ceg_net566), .I1(n9879), .O(ceg_net1361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__13853.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__13854 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(n9856), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n899 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__13854.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__13855 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .O(n9902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__13855.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__13856 (.I0(n9854), .I1(n9876), .I2(n9902), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n898 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__13856.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__13857 (.I0(n9851), .I1(n9868), .O(ceg_net616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__13857.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__13858 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] ), 
            .I2(n9852), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__13858.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__13859 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] ), 
            .I3(n9852), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n844 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__13859.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__13860 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3] ), 
            .O(n9903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h807f */ ;
    defparam LUT__13860.LUTMASK = 16'h807f;
    EFX_LUT4 LUT__13861 (.I0(n9903), .I1(n9852), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13861.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13862 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3] ), 
            .O(n9904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13862.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13863 (.I0(n9904), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] ), 
            .I2(n9852), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n842 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__13863.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__13864 (.I0(n9904), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] ), 
            .O(n9905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13864.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13865 (.I0(n9905), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] ), 
            .I2(n9852), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n841 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__13865.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__13866 (.I0(n9905), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6] ), 
            .I3(n9852), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n840 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__13866.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__13867 (.I0(n9904), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6] ), 
            .O(n9906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13867.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13868 (.I0(n9906), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .I2(n9852), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n839 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__13868.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__13883 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] ), 
            .I2(n9853), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__13883.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__13884 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2] ), 
            .I3(n9853), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n850 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__13884.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__13885 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n869 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13885.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13886 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n868 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13886.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13887 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n867 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13887.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13888 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n866 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13888.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13889 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n865 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13889.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13890 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n864 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13890.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13891 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n863 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13891.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13892 (.I0(n9854), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0] ), 
            .O(n9913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13892.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13893 (.I0(n9854), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1] ), 
            .I3(n9884), .O(n9914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__13893.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__13894 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n9915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7e7 */ ;
    defparam LUT__13894.LUTMASK = 16'he7e7;
    EFX_LUT4 LUT__13895 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] ), 
            .I2(n9885), .I3(n9866), .O(n9916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__13895.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__13896 (.I0(n9915), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] ), 
            .I2(n9916), .O(n9917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__13896.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__13897 (.I0(n9913), .I1(n9914), .I2(n9868), .I3(n9917), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n878 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0ff */ ;
    defparam LUT__13897.LUTMASK = 16'hb0ff;
    EFX_LUT4 LUT__13898 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] ), 
            .I2(n9885), .O(n9918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__13898.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__13899 (.I0(n9854), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2] ), 
            .I3(n9884), .O(n9919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__13899.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__13900 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(n9918), .I2(n9919), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n9920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__13900.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__13901 (.I0(n9920), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I2(n9915), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n877 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f11 */ ;
    defparam LUT__13901.LUTMASK = 16'h1f11;
    EFX_LUT4 LUT__13902 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] ), 
            .I2(n9885), .O(n9921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__13902.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__13903 (.I0(n9854), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3] ), 
            .I3(n9884), .O(n9922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__13903.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__13904 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(n9921), .I2(n9922), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n9923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__13904.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__13905 (.I0(n9923), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I2(n9915), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n876 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f11 */ ;
    defparam LUT__13905.LUTMASK = 16'h1f11;
    EFX_LUT4 LUT__13906 (.I0(n9854), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4] ), 
            .I3(n9884), .O(n9924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__13906.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__13907 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] ), 
            .I2(n9885), .I3(n9866), .O(n9925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__13907.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__13908 (.I0(n9915), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] ), 
            .I2(n9925), .O(n9926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__13908.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__13909 (.I0(n9913), .I1(n9924), .I2(n9868), .I3(n9926), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n875 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0ff */ ;
    defparam LUT__13909.LUTMASK = 16'hb0ff;
    EFX_LUT4 LUT__13910 (.I0(n9854), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5] ), 
            .I3(n9884), .O(n9927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__13910.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__13911 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] ), 
            .I2(n9885), .I3(n9866), .O(n9928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__13911.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__13912 (.I0(n9913), .I1(n9927), .I2(n9868), .I3(n9928), 
            .O(n9929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__13912.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__13913 (.I0(n9915), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] ), 
            .I2(n9929), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n874 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__13913.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__13914 (.I0(n9854), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6] ), 
            .I3(n9884), .O(n9930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__13914.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__13915 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] ), 
            .I2(n9885), .I3(n9866), .O(n9931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__13915.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__13916 (.I0(n9915), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] ), 
            .I2(n9931), .O(n9932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__13916.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__13917 (.I0(n9913), .I1(n9930), .I2(n9868), .I3(n9932), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n873 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0ff */ ;
    defparam LUT__13917.LUTMASK = 16'hb0ff;
    EFX_LUT4 LUT__13918 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] ), 
            .I2(n9885), .O(n9933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__13918.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__13919 (.I0(n9854), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7] ), 
            .I3(n9884), .O(n9934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__13919.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__13920 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(n9933), .I2(n9934), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n9935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__13920.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__13921 (.I0(n9935), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I2(n9915), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n872 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f11 */ ;
    defparam LUT__13921.LUTMASK = 16'h1f11;
    EFX_LUT4 LUT__13929 (.I0(oAdv7511SdaOe), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(iAdv7511Sda), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n9936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3 */ ;
    defparam LUT__13929.LUTMASK = 16'hedf3;
    EFX_LUT4 LUT__13930 (.I0(n9876), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I2(n9936), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n9937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__13930.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__13931 (.I0(n9937), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n828 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13931.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13932 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I1(n9875), .I2(n9872), .I3(n9878), .O(n9938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__13932.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__13933 (.I0(n9849), .I1(n9868), .I2(n9938), .O(ceg_net1471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__13933.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__13934 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I2(n9864), .O(n9939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__13934.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__13935 (.I0(n9939), .I1(n9849), .I2(n9896), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n9940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__13935.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__13936 (.I0(n9940), .I1(n9856), .I2(n9893), .I3(n9869), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n827 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888 */ ;
    defparam LUT__13936.LUTMASK = 16'hf888;
    EFX_LUT4 LUT__13937 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I1(n9849), .I2(n9866), .I3(n9938), .O(n9941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__13937.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__13938 (.I0(n9868), .I1(n9895), .I2(n9941), .O(ceg_net1480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f8f */ ;
    defparam LUT__13938.LUTMASK = 16'h8f8f;
    EFX_LUT4 LUT__13939 (.I0(n9876), .I1(n9892), .I2(n9939), .I3(n9856), 
            .O(n9942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__13939.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__13940 (.I0(n9869), .I1(n9888), .I2(n9942), .I3(n9871), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n826 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__13940.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__13941 (.I0(n9857), .I1(n9849), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n9943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8cf */ ;
    defparam LUT__13941.LUTMASK = 16'hf8cf;
    EFX_LUT4 LUT__13942 (.I0(n9943), .I1(n9856), .I2(n9938), .O(ceg_net1488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__13942.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__13943 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[0] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[1] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[3] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rVpos[4] ), .O(n9944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13943.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13944 (.I0(n9944), .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[5] ), 
            .O(n9945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13944.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13945 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[5] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[3] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[4] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rVpos[2] ), .O(n9946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__13945.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__13946 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[7] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[8] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[9] ), 
            .O(n9947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__13946.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__13947 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[11] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[6] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[10] ), 
            .I3(n9947), .O(n9948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__13947.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__13948 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[2] ), 
            .I1(n9945), .I2(n9946), .I3(n9948), .O(\MVideoPostProcess/mVideoTimingGen/qVrange )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__13948.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__13949 (.I0(\MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n251 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__13949.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__13950 (.I0(\MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] ), 
            .O(n9949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__13950.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__13951 (.I0(n9949), .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n250 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13951.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13952 (.I0(\MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] ), 
            .O(n9950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13952.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13953 (.I0(n9950), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n249 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__13953.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__13954 (.I0(n9950), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] ), 
            .O(n9951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13954.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13955 (.I0(n9951), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__13955.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__13956 (.I0(n9951), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] ), 
            .O(n9952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13956.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13957 (.I0(n9952), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n247 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__13957.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__13958 (.I0(n9952), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n246 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__13958.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__13959 (.I0(n9952), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] ), .O(n9953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13959.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13960 (.I0(n9953), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n245 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__13960.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__13961 (.I0(n9953), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n244 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__13961.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__13962 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n700 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13962.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13963 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n705 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13963.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13964 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n710 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__13964.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__13965 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3] ), 
            .O(n9954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13965.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13966 (.I0(n9954), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n715 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13966.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13967 (.I0(n9954), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n720 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13967.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13968 (.I0(n9954), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n725 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__13968.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__13969 (.I0(n9954), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6] ), 
            .O(n9955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13969.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13970 (.I0(n9955), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n730 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13970.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13971 (.I0(n9955), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7] ), 
            .O(n9956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13971.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13972 (.I0(n9956), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n735 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13972.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13973 (.I0(n9956), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n740 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13973.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13974 (.I0(n9956), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9] ), 
            .O(n9957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13974.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13975 (.I0(n9957), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n745 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13975.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13976 (.I0(n9957), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n750 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13976.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13977 (.I0(n9957), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n755 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__13977.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__13978 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] ), 
            .O(n9958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13978.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13979 (.I0(n9956), .I1(n9958), .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9] ), 
            .O(n9959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13979.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13980 (.I0(n9959), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n760 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13980.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13981 (.I0(n9959), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n765 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13981.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13982 (.I0(n9959), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__13982.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__13983 (.I0(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] ), .O(\MVideoPostProcess/inst_adv7511_config/n780 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13983.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13984 (.I0(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n785 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13984.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13985 (.I0(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3] ), .O(\MVideoPostProcess/inst_adv7511_config/n790 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__13985.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__13986 (.I0(n9845), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n795 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13986.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13987 (.I0(n9845), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] ), .O(\MVideoPostProcess/inst_adv7511_config/n800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13987.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13988 (.I0(n9845), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n805 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__13988.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__13989 (.I0(n9846), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13989.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13990 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n276 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__13990.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__13991 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n275 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__13991.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__13992 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[3] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n274 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__13992.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__13993 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n273 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__13993.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__13994 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n272 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__13994.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__13995 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[6] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n271 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__13995.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__13996 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[7] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__13996.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__13997 (.I0(n9948), .I1(n9945), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[2] ), 
            .O(n9960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13997.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13998 (.I0(n9960), .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[0] ), 
            .O(\MVideoPostProcess/mVideoTimingGen/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13998.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13999 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[3] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[5] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[6] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rHpos[8] ), .O(n9961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13999.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__14000 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[9] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[10] ), .I2(n9961), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rHpos[11] ), .O(n9962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__14000.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__14001 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[0] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[1] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[2] ), 
            .O(n9675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14001.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14002 (.I0(n9962), .I1(n9675), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[4] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rHpos[7] ), .O(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__14002.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__14003 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[4] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[5] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[3] ), 
            .I3(n9947), .O(n9963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__14003.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__14004 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[7] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[8] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[9] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rHpos[10] ), .O(n9964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14004.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14005 (.I0(n9964), .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[11] ), 
            .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[11] ), .O(n9965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__14005.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__14006 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[6] ), 
            .I1(n9963), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[10] ), 
            .I3(n9965), .O(\MVideoPostProcess/mVideoTimingGen/qVde )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__14006.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__14007 (.I0(\MVideoPostProcess/rVtgRST[2] ), .I1(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
            .O(\MVideoPostProcess/mVideoTimingGen/n267 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__14007.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__14008 (.I0(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3 ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/dff_11/i4_pre ), .O(\MVideoPostProcess/mVideoTimingGen/rHSync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14008.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14009 (.I0(n9960), .I1(n492), .O(\MVideoPostProcess/mVideoTimingGen/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14009.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14010 (.I0(n9960), .I1(n3699), .O(\MVideoPostProcess/mVideoTimingGen/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14010.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14011 (.I0(n9960), .I1(n3693), .O(\MVideoPostProcess/mVideoTimingGen/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14011.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14012 (.I0(n9960), .I1(n3691), .O(\MVideoPostProcess/mVideoTimingGen/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14012.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14013 (.I0(n9960), .I1(n3683), .O(\MVideoPostProcess/mVideoTimingGen/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14013.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14014 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[3] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[4] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[5] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rHpos[11] ), .O(n9966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__14014.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__14015 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[2] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[4] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[7] ), 
            .I3(n9962), .O(n9967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__14015.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__14016 (.I0(n9966), .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[6] ), 
            .I2(n9964), .I3(n9967), .O(\MVideoPostProcess/mVideoTimingGen/qHrange )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff80 */ ;
    defparam LUT__14016.LUTMASK = 16'hff80;
    EFX_LUT4 LUT__14017 (.I0(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_pre ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3 ), .O(\MVideoPostProcess/mVideoTimingGen/rVSync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14017.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14018 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .O(n9968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14018.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14019 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n9969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14019.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14020 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n9970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14020.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14021 (.I0(n9969), .I1(n9970), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n9971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001 */ ;
    defparam LUT__14021.LUTMASK = 16'h1001;
    EFX_LUT4 LUT__14022 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(n9972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb00b */ ;
    defparam LUT__14022.LUTMASK = 16'hb00b;
    EFX_LUT4 LUT__14023 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n9973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14023.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14024 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n9974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb00b */ ;
    defparam LUT__14024.LUTMASK = 16'hb00b;
    EFX_LUT4 LUT__14025 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n9975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14025.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14026 (.I0(n9972), .I1(n9973), .I2(n9974), .I3(n9975), 
            .O(n9976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14026.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14027 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(n9971), .I3(n9976), .O(n9977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14027.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14028 (.I0(n9977), .I1(n9968), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14028.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14029 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(n9978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14029.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14030 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n9979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14030.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14031 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n9980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14031.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14032 (.I0(n9979), .I1(n9980), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n9981)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14032.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14033 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n9982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__14033.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__14034 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
            .I1(n9982), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n9983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__14034.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__14035 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n9984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__14035.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__14036 (.I0(n9981), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(n9983), .I3(n9984), .O(n9985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__14036.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__14037 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n9986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__14037.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__14038 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n9987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14038.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14039 (.I0(n9987), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(n9988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14039.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14040 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] ), 
            .I1(n9986), .I2(n9988), .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n9989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__14040.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__14041 (.I0(n9979), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(n9990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14041.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14042 (.I0(n9969), .I1(n9990), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .O(n9991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be */ ;
    defparam LUT__14042.LUTMASK = 16'he7be;
    EFX_LUT4 LUT__14043 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n9992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__14043.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__14044 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n9993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14044.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14045 (.I0(n9987), .I1(n9993), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n9994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14045.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14046 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] ), 
            .I1(n9992), .I2(n9994), .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n9995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__14046.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__14047 (.I0(n9989), .I1(n9991), .I2(n9995), .O(n9996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__14047.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__14048 (.I0(n9979), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .O(n9997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14048.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14049 (.I0(n9970), .I1(n9997), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n9998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be */ ;
    defparam LUT__14049.LUTMASK = 16'he7be;
    EFX_LUT4 LUT__14050 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] ), 
            .I1(n9986), .I2(n9987), .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n9999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__14050.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__14051 (.I0(n9982), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7e7 */ ;
    defparam LUT__14051.LUTMASK = 16'he7e7;
    EFX_LUT4 LUT__14052 (.I0(n9999), .I1(n10000), .I2(n9981), .I3(n9984), 
            .O(n10001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110 */ ;
    defparam LUT__14052.LUTMASK = 16'h0110;
    EFX_LUT4 LUT__14053 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .O(n10002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__14053.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__14054 (.I0(n10002), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I3(n9978), .O(n10003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__14054.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__14055 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb00b */ ;
    defparam LUT__14055.LUTMASK = 16'hb00b;
    EFX_LUT4 LUT__14056 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I3(n10004), .O(n10005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100 */ ;
    defparam LUT__14056.LUTMASK = 16'h7100;
    EFX_LUT4 LUT__14057 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .O(n10006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14057.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14058 (.I0(n9980), .I1(n9992), .I2(n10006), .I3(n9979), 
            .O(n10007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9ff3 */ ;
    defparam LUT__14058.LUTMASK = 16'h9ff3;
    EFX_LUT4 LUT__14059 (.I0(n10005), .I1(n10003), .I2(n10007), .O(n10008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__14059.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__14060 (.I0(n10005), .I1(n10003), .I2(n9971), .I3(n9976), 
            .O(n10009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__14060.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__14061 (.I0(n9998), .I1(n10008), .I2(n10001), .I3(n10009), 
            .O(n10010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__14061.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__14062 (.I0(n9985), .I1(n9996), .I2(n9978), .I3(n10010), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qFullAllmost )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h80ff */ ;
    defparam LUT__14062.LUTMASK = 16'h80ff;
    EFX_LUT4 LUT__14063 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14063.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14064 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n483 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14064.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14065 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n488 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14065.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14066 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(n10011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14066.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14067 (.I0(n10011), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n493 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14067.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14068 (.I0(n10011), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14068.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14069 (.I0(n9987), .I1(n10011), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n503 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14069.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14070 (.I0(n9987), .I1(n10011), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n508 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14070.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14071 (.I0(n9979), .I1(n10011), .O(n10012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14071.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14072 (.I0(n10012), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n513 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14072.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14073 (.I0(n9997), .I1(n10011), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n518 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14073.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14074 (.I0(n10012), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n523 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14074.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14075 (.I0(n10012), .I1(n9980), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n528 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14075.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14076 (.I0(n9981), .I1(n10011), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n533 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14076.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14077 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14077.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14078 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14078.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14079 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14079.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14080 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14080.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14081 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14081.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14082 (.I0(n10014), .I1(n10015), .I2(n10016), .I3(n10017), 
            .O(n10018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14082.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14083 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14083.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14084 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(n10018), .I3(n10019), .O(n10020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14084.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14085 (.I0(n10020), .I1(n10013), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14085.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14086 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14086.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14087 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14087.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14088 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14088.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14089 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14089.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14090 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14090.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14091 (.I0(n10022), .I1(n10023), .I2(n10024), .I3(n10025), 
            .O(n10026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14091.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14092 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14092.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14093 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(n10026), .I3(n10027), .O(n10028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14093.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14094 (.I0(n10028), .I1(n10021), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14094.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14095 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14095.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14096 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n10030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14096.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14097 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14097.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14098 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14098.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14099 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14099.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14100 (.I0(n10030), .I1(n10031), .I2(n10032), .I3(n10033), 
            .O(n10034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14100.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14101 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14101.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14102 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(n10034), .I3(n10035), .O(n10036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14102.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14103 (.I0(n10036), .I1(n10029), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14103.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14104 (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14104.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14105 (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14105.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14106 (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14106.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14107 (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14107.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14108 (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14108.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14109 (.I0(n10038), .I1(n10039), .I2(n10040), .I3(n10041), 
            .O(n10042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14109.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14110 (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14110.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14111 (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(n10042), .I3(n10043), .O(n10044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14111.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14112 (.I0(n10044), .I1(n10037), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14112.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14113 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14113.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14114 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14114.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14115 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14115.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14116 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14116.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14117 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14117.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14118 (.I0(n10046), .I1(n10047), .I2(n10048), .I3(n10049), 
            .O(n10050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14118.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14119 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14119.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14120 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0] ), 
            .I2(n10050), .I3(n10051), .O(n10052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14120.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14121 (.I0(n10052), .I1(n10045), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14121.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14122 (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14122.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14123 (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .I2(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14123.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14124 (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14124.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14125 (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14125.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14126 (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14126.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14127 (.I0(n10054), .I1(n10055), .I2(n10056), .I3(n10057), 
            .O(n10058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14127.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14128 (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14128.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14129 (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(n10058), .I3(n10059), .O(n10060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14129.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14130 (.I0(n10060), .I1(n10053), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14130.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14131 (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14131.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14132 (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14132.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14133 (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .I2(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14133.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14134 (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n10064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14134.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14135 (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14135.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14136 (.I0(n10062), .I1(n10063), .I2(n10064), .I3(n10065), 
            .O(n10066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14136.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14137 (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14137.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14138 (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0] ), 
            .I2(n10066), .I3(n10067), .O(n10068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14138.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14139 (.I0(n10068), .I1(n10061), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14139.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14140 (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14140.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14141 (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14141.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14142 (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14142.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14143 (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14143.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14144 (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14144.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14145 (.I0(n10070), .I1(n10071), .I2(n10072), .I3(n10073), 
            .O(n10074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14145.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14146 (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14146.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14147 (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(n10074), .I3(n10075), .O(n10076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14147.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14148 (.I0(n10076), .I1(n10069), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14148.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14149 (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14149.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14150 (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14150.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14151 (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14151.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14152 (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(n10080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14152.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14153 (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14153.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14154 (.I0(n10078), .I1(n10079), .I2(n10080), .I3(n10081), 
            .O(n10082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14154.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14155 (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14155.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14156 (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0] ), 
            .I2(n10082), .I3(n10083), .O(n10084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14156.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14157 (.I0(n10084), .I1(n10077), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14157.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14158 (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14158.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14159 (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14159.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14160 (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14160.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14161 (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14161.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14162 (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14162.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14163 (.I0(n10086), .I1(n10087), .I2(n10088), .I3(n10089), 
            .O(n10090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14163.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14164 (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14164.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14165 (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(n10090), .I3(n10091), .O(n10092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14165.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14166 (.I0(n10092), .I1(n10085), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14166.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14167 (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14167.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14168 (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14168.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14169 (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14169.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14170 (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(n10096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14170.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14171 (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14171.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14172 (.I0(n10094), .I1(n10095), .I2(n10096), .I3(n10097), 
            .O(n10098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14172.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14173 (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14173.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14174 (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0] ), 
            .I2(n10098), .I3(n10099), .O(n10100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14174.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14175 (.I0(n10100), .I1(n10093), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14175.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14176 (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14176.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14177 (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14177.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14178 (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14178.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14179 (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14179.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14180 (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14180.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14181 (.I0(n10102), .I1(n10103), .I2(n10104), .I3(n10105), 
            .O(n10106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14181.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14182 (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14182.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14183 (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(n10106), .I3(n10107), .O(n10108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14183.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14184 (.I0(n10108), .I1(n10101), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14184.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14185 (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14185.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14186 (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(n10110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14186.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14187 (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14187.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14188 (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14188.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14189 (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14189.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14190 (.I0(n10110), .I1(n10111), .I2(n10112), .I3(n10113), 
            .O(n10114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14190.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14191 (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14191.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14192 (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(n10114), .I3(n10115), .O(n10116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14192.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14193 (.I0(n10116), .I1(n10109), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14193.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14194 (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14194.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14195 (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14195.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14196 (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14196.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14197 (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14197.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14198 (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .I2(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14198.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14199 (.I0(n10118), .I1(n10119), .I2(n10120), .I3(n10121), 
            .O(n10122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14199.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14200 (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14200.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14201 (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(n10122), .I3(n10123), .O(n10124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14201.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14202 (.I0(n10124), .I1(n10117), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14202.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14203 (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14203.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14204 (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14204.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14205 (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14205.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14206 (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14206.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14207 (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .I2(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14207.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14208 (.I0(n10126), .I1(n10127), .I2(n10128), .I3(n10129), 
            .O(n10130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14208.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14209 (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14209.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14210 (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(n10130), .I3(n10131), .O(n10132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14210.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14211 (.I0(n10132), .I1(n10125), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14211.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14212 (.I0(\genblk1.genblk1[0].mPulseGenerator/rSft[2] ), 
            .I1(\genblk1.genblk1[0].mPulseGenerator/rSft[1] ), .I2(\genblk1.genblk1[0].mPulseGenerator/rSft[0] ), 
            .O(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf */ ;
    defparam LUT__14212.LUTMASK = 16'hbfbf;
    EFX_LUT4 LUT__14213 (.I0(n3370), .I1(n3368), .I2(n3366), .I3(n3364), 
            .O(n10133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__14213.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__14214 (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[3] ), 
            .I1(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[4] ), .I2(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_0_q ), 
            .O(n10134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14214.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14215 (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] ), 
            .I1(n1219), .I2(n1193), .O(n9476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__14215.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__14216 (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[10] ), 
            .I1(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[11] ), .I2(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[9] ), 
            .I3(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[12] ), .O(n10135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__14216.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__14217 (.I0(n10134), .I1(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_1_q ), 
            .I2(n10135), .O(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f7f */ ;
    defparam LUT__14217.LUTMASK = 16'h7f7f;
    EFX_LUT4 LUT__14218 (.I0(\genblk1.genblk1[3].mPulseGenerator/rSft[2] ), 
            .I1(\genblk1.genblk1[3].mPulseGenerator/rSft[1] ), .I2(\genblk1.genblk1[3].mPulseGenerator/rSft[0] ), 
            .O(\genblk1.genblk1[3].mPulseGenerator/equal_6/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf */ ;
    defparam LUT__14218.LUTMASK = 16'hbfbf;
    EFX_LUT4 LUT__14219 (.I0(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[0] ), 
            .I1(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] ), .O(\genblk1.genblk1[3].mPulseGenerator/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14219.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14220 (.I0(\genblk1.genblk1[4].mPulseGenerator/rSft[2] ), 
            .I1(\genblk1.genblk1[4].mPulseGenerator/rSft[1] ), .I2(\genblk1.genblk1[4].mPulseGenerator/rSft[0] ), 
            .O(\genblk1.genblk1[4].mPulseGenerator/equal_6/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf */ ;
    defparam LUT__14220.LUTMASK = 16'hbfbf;
    EFX_LUT4 LUT__14221 (.I0(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[0] ), 
            .I1(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] ), .O(\genblk1.genblk1[4].mPulseGenerator/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14221.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14222 (.I0(\la0_probe3[0] ), .I1(\la0_probe3[1] ), .O(la0_probe1)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14222.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13628 (.I0(pll_inst1_LOCKED), .I1(pll_inst2_LOCKED), .O(oLed[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13628.LUTMASK = 16'h8888;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_1  (.D(n9476), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_1_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, INIT_VALUE=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_1 .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_1 .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_1 .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_1 .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_1 .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_1 .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_1 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_0  (.D(n10133), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n25 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_0_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, INIT_VALUE=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_0 .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_0 .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_0 .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_0 .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_0 .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_0 .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_0 .SR_SYNC_PRIORITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_FF_cc8bc306_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_cc8bc306_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_cc8bc306_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__10_10_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__10_10_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__16_16_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__8_8_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_SRL8_cc8bc306_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__1_1_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_cc8bc306__2_2_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_173
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_174
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_175
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_176
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_177
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_178
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_179
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_180
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_181
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_182
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_183
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_184
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_185
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_186
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_187
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_188
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_189
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_190
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_191
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_192
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_193
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_194
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_195
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_196
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_197
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_198
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_199
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_200
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_201
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_202
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_203
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_204
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_205
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_206
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_207
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_208
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_209
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_210
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_211
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_212
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_213
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_214
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_cc8bc306_215
// module not written out since it is a black box. 
//

