module SEG10_COUNT_sim;

endmodule