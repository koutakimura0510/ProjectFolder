//----------------------------------------------------------
// Create 2022/02/05
// Author koutakimura
// -
// FIFOコントロールモジュール
// この回路を使用する上位モジュールでは下記の内容でデータのやり取りを行う
// 1.書き込み時はoFullのみ確認すれば良い
// 2.読み込み時はoEMPとoRdVを確認すれば良い
//
// 2022/02/26
// 処理の流れが分かりにくいため、全体をパイプライン処理に更新
// RE Active時 3CLK後に RVD Assert データが出力される
// 
// 2022/03/13
// 動作周波数を上げるため全体構成見直し、パイプライン処理中止
//
// 2022-03-21
// ReadEnableから 2レイテンシでデータ出力する構造に変更、ユーザが意識せずともハンドシェイクが上手く行く用に変更
//
// 2022-09-06
// コーディング規則に則りソースコードの修正
// 
//----------------------------------------------------------
module fifoController #(
    parameter 					pFifoDepth        	= 1024,		// FIFO BRAMのサイズ指定
    parameter 					pFifoBitWidth     	= 8,		// bitサイズ
	parameter 					pFifoCascade		= 1,     	// BRAM使用個数
	parameter					pFullAlMost 		= 6,		// 指定値、早く full 出力
	parameter	[0:0]			pFullRst 			= 1'b0,
	parameter	[0:0]			pEmpRst 			= 1'b1,
	parameter					pFifoBlockRam		= "yes",	// yes BRAM, no reg
	parameter					pAddrWidth			= fBitWidth(pFifoDepth)
)(
	// src side
    input   [pFifoBitWidth-1:0] iWd,        // write data
    input                       iWe,        // write enable Active High
    output                      oFull,      // Fifo Full Assert, Active High
	// dst side
    output  [pFifoBitWidth-1:0] oRd,        // read data
    input                       iRe,        // read enable Active High
    output                      oRvd,       // Valid Data
    output                      oEmp,       // Fifo Empty
	//
    input                       iRST,
    input                       iCLK
);
	// .iWd	(),				.iWe	(),
	// .oFull	(),
	// .oRd	(),				.iRe	(),
	// .oRvd	(),				.oEmp	(),
	// .iRST	(qSRST),		.iCLK	(iSCLK)


//-----------------------------------------------------------------------------
// アドレスの更新
//-----------------------------------------------------------------------------
reg [pAddrWidth-1:0] rWa, rRa, rRaOld;
reg qWe, qRe;

always @(posedge iCLK)
begin
    if (iRST)       rWa <= {pAddrWidth{1'b0}};
    else if (qWe)   rWa <= rWa + 1'b1;
    else            rWa <= rWa;
	//
    if (iRST)      	rRa <= {pAddrWidth{1'b0}};
    else if (qRe)  	rRa <= rRa + 1'b1;
    else           	rRa <= rRa;
	// 前回のrpが更新されていたら新規データを出力できる状態と判断する
    if (iRST)   	rRaOld <= {pAddrWidth{1'b0}};
    else        	rRaOld <= rRa;
end


//----------------------------------------------------------
// ハンドシェイク信号出力
//----------------------------------------------------------
localparam lpFullAlMost = pFullAlMost + 1;

reg 					rFull;						assign oFull = rFull;
reg 					rEmp;						assign oEmp  = rEmp;
reg 					rRvd;						assign oRvd  = rRvd;
reg 					qFullAllmost, qEmp, qRvd;
reg [pFullAlMost-1:0] 	qFull;
reg [pAddrWidth-1:0] 	qWAn [0:pFullAlMost];

always @(posedge iCLK)
begin
	if (iRST)				rFull <= pFullRst;
	else if (qFullAllmost)	rFull <= 1'b1;
	else					rFull <= 1'b0;

	if (iRST)				rEmp <= pEmpRst;
	else if (qEmp)			rEmp <= 1'b1;
	else					rEmp <= 1'b0;

	if (iRST)				rRvd <= 1'b0;
	else if	(qRvd)			rRvd <= 1'b1;
	else					rRvd <= 1'b0;
end
//
integer n;

generate
	always @*
	begin
		for (n = 1; n < lpFullAlMost; n = n + 1)
		begin
			qWAn[n-1]   <= rWa + n;
			qFull[n-1]	<= (qWAn[n-1] == rRa);
		end
		qFullAllmost <= |{qFull};
	end
endgenerate

always @*
begin
    qEmp <= (rWa == rRa);
    qRvd <= (rRa != rRaOld);
    qWe  <= iWe;
    qRe  <= iRe & (~qEmp);
end


//----------------------------------------------------------
// FIFO 動作
//----------------------------------------------------------
wire	[pFifoBitWidth-1:0] wRd;					assign oRd = wRd;

genvar m;

generate
	for (m = 0; m < pFifoCascade; m = m + 1)
	begin
		userFifo #(
			.pBuffDepth    	(pFifoDepth),
			.pBitWidth     	(pFifoBitWidth),
			.pAddrWidth    	(pAddrWidth),
			.pFifoBlockRam	(pFifoBlockRam)
		) USER_FIFO (
			// write
			.iWD(iWd[(m+1)*(pFifoBitWidth/pFifoCascade)-1:m*(pFifoBitWidth/pFifoCascade)]),
			.iWA(rWa),			.iWE(qWe),
			// read
			.oRD(wRd[(m+1)*(pFifoBitWidth/pFifoCascade)-1:m*(pFifoBitWidth/pFifoCascade)]),
			.iRA(rRa),
			.iClk(iCLK)
		);
	end
endgenerate


//-----------------------------------------------------------------------------
// msb側の1を検出しbit幅を取得する
//-----------------------------------------------------------------------------
function[  7:0]	fBitWidth;
    input [31:0] iVAL;
    integer			i;

    begin
    // fBitWidth = 1;
        for (i = 0; i < 32; i = i+1 )
        begin
            if (iVAL[i]) 
            begin
                fBitWidth = i+1;
            end
        end

        if (fBitWidth != 1)
        begin
            fBitWidth = fBitWidth - 1;
        end
    end
endfunction
////////////////////////////////////////////////////////////
endmodule