//-----------------------------------------------------------------------------
// Create  2023/1/7
// Author  kimura
// Editor  VSCode ver1.70.0
// -
// Dual Port RAM のプリミティブをインスタンスする
// 
//-----------------------------------------------------------------------------
module EfxRam10Primitive #(
    parameter 					pBitWidth  		= 16,	// Data Width
    parameter 					pAddrWidth 		= 13
)(
	// Write Side
    input	[pBitWidth-1:0]		iWd,    // write data
    input	[pAddrWidth-1:0]	iWa,    // write addr
    input						iWe,    // write enable
	// Read Side
    output	[pBitWidth-1:0]		oRd,    // read data
    input	[pAddrWidth-1:0]	iRa,    // read address
	input 						iRe,
	// common
	input 						iRST,
    input						iCLK
);

generate
	if (pAddrWidth == 13)
	begin
		EFX_RAM10 # (
			.WCLK_POLARITY(1'b1), 		// wclk 	polarity
			.WCLKE_POLARITY(1'b1), 		// wclke 	polarity
			.WADDREN_POLARITY(1'b1), 	// waddren 	polarity
			.WE_POLARITY(2'b11), 		// we 		polarity
			.RCLK_POLARITY(1'b1), 		// rclk 	polarity
			.RE_POLARITY(1'b1), 		// re 		polarity
			.RST_POLARITY(1'b1), 		// rst 		polarity
			.RADDREN_POLARITY(1'b1), 	// raddren 	polarity
			.READ_WIDTH(pBitWidth),		// read 	width
			.WRITE_WIDTH(pBitWidth),	// write 	width
			.OUTPUT_REG(1'b1), 			// Output 	register enable
			.WRITE_MODE("READ_FIRST"), 	// write 	mode
			.RESET_RAM("ASYNC"), 		// reset 	mode on ram
			.RESET_OUTREG("ASYNC"), 	// reset 	mode on output register
			// 256-bit INIT string
			.INIT_0 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_1 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_2 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_3 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_4 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_5 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_6 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_7 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_8 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_9 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_A (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_B (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_C (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_D (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_E (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_F (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_10 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_11 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_12 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_13 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_14 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_15 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_16 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_17 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_18 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_19 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_1A (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_1B (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_1C (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_1D (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_1E (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_1F (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_20 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_21 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_22 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_23 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_24 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_25 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_26 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_27 (256'h0000000000000000000000000000000000000000000000000000000000000000)
		)
		ram10_inst (
			.WCLK(iCLK), 		// write clk
			.WE({2{iWe}}),		// 2-bit write enable, [1]=[15:8], [0]=[7:0]
			.WCLKE(1'b1), 		// write clk enable
			.WADDREN(iWe),	 	// write address enable
			.WDATA(iWd), 		// write data input
			.WADDR(iWa), 		// write address input
			.RCLK(iCLK), 		// read clk
			.RE(iRe), 			// read enable
			.RST(iRST),			// reset
			.RADDREN(iRe),	 	// read address enable
			.RDATA(oRd), 		// read data output
			.RADDR(iRa) 		// read address input
		);
	end
	else
	begin
		EFX_RAM10 # (
			.WCLK_POLARITY(1'b1), 		// wclk 	polarity
			.WCLKE_POLARITY(1'b1), 		// wclke 	polarity
			.WADDREN_POLARITY(1'b1), 	// waddren 	polarity
			.WE_POLARITY(2'b11), 		// we 		polarity
			.RCLK_POLARITY(1'b1), 		// rclk 	polarity
			.RE_POLARITY(1'b1), 		// re 		polarity
			.RST_POLARITY(1'b1), 		// rst 		polarity
			.RADDREN_POLARITY(1'b1), 	// raddren 	polarity
			.READ_WIDTH(pBitWidth),		// read 	width
			.WRITE_WIDTH(pBitWidth),	// write 	width
			.OUTPUT_REG(1'b1), 			// Output 	register enable
			.WRITE_MODE("READ_FIRST"), 	// write 	mode
			.RESET_RAM("ASYNC"), 		// reset 	mode on ram
			.RESET_OUTREG("ASYNC"), 	// reset 	mode on output register
			// 256-bit INIT string
			.INIT_0 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_1 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_2 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_3 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_4 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_5 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_6 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_7 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_8 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_9 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_A (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_B (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_C (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_D (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_E (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_F (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_10 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_11 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_12 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_13 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_14 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_15 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_16 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_17 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_18 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_19 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_1A (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_1B (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_1C (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_1D (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_1E (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_1F (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_20 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_21 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_22 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_23 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_24 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_25 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_26 (256'h0000000000000000000000000000000000000000000000000000000000000000),
			.INIT_27 (256'h0000000000000000000000000000000000000000000000000000000000000000)
		)
		ram10_inst (
			.WCLK(iCLK), 		// write clk
			.WE({2{iWe}}),		// 2-bit write enable, [1]=[15:8], [0]=[7:0]
			.WCLKE(1'b1), 		// write clk enable
			.WADDREN(iWe),	 	// write address enable
			.WDATA(iWd), 		// write data input
			.WADDR({{(13-pAddrWidth){1'b0}},iWa}), // write address input
			.RCLK(iCLK), 		// read clk
			.RE(iRe), 			// read enable
			.RST(iRST),			// reset
			.RADDREN(iRe),	 	// read address enable
			.RDATA(oRd), 		// read data output
			.RADDR({{(13-pAddrWidth){1'b0}},iRa}) // read address input
		);
	end
endgenerate

endmodule
