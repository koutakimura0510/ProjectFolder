//----------------------------------------------------------
// Create 2022/08/31
// Author koutakimura
// -
// 指定範囲で指定色の四角形データを出力する
// 
// 2022-09-29 座標が画面外の場合のドットデータ生成に対応
// 
//----------------------------------------------------------
module DotSquareGen #(
	parameter	pVHAW  = 11,
	parameter	pVVAW  = 11,
	parameter	pColorDepth = 16
)(
	// Pixel Output
	output	[pColorDepth-1:0]	oPd,		// Pixel Data
	output 						oPv,		// Pixel Valid
	// Control Status
	input	[pColorDepth-1:0]	iColor,		// 描画色
	input	[pVHAW-1:0]	iHpos,				// 現在の横幅の座標
	input	[pVVAW-1:0]	iVpos,				// 現在の立幅の座標
	input signed	[pVHAW:0]	iDLeftX,	// 描画開始 X座標 Draw X Start
	input signed	[pVHAW:0]	iDRightX,	// 描画終了 X座標 Draw X End
	input signed	[pVVAW:0]	iDTopY,		// 描画開始 Y座標 Draw Y Start
	input signed	[pVVAW:0]	iDUnderY,	// 描画終了 Y座標 Draw Y End
	// Common
	input	iRST,
	input	iCLK
);


//-----------------------------------------------------------------------------
// 符号拡張
//-----------------------------------------------------------------------------
wire signed [pVHAW:0] wHpos = {1'b0, iHpos};
wire signed [pVVAW:0] wVpos = {1'b0, iVpos};


//-----------------------------------------------------------------------------
// 指定色のデータ及び範囲外であれば透過値最大のデータを出力
// 画面外に座標データがはみ出ても、範囲内のドットデータは描画するようにする
//-----------------------------------------------------------------------------
reg [pColorDepth-1:0] rPd;		assign oPd = qCke ? iColor : 0; //rPd;
reg rPv;						assign oPv = rPv;
reg qCke;
reg [3:0] qPosMatch;

always @(posedge iCLK)
begin
	if (qCke) 		rPd <= iColor;
    else 			rPd <= {pColorDepth{1'b0}};
	
	if (iRST) 		rPv <= 1'b0;
	else 			rPv <= qCke;
end

always @*
begin
	qPosMatch[0] <= (iDLeftX <= wHpos);
	qPosMatch[1] <= (wHpos 	 <  iDRightX);
	qPosMatch[2] <= (iDTopY  <= wVpos);
	qPosMatch[3] <= (wVpos   <  iDUnderY);
	qCke 		 <= &(qPosMatch);
end

endmodule