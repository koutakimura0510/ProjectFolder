//////////////////////////////////////////////////////////////////////////////////////////
//           _____       
//          / _______    Copyright (C) 2013-2022 Efinix Inc. All rights reserved.
//         / /       \   
//        / /  ..    /   
//       / / .'     /    
//    __/ /.'      /     Description:
//   __   \       /      Top IP Module = efx_csi2_tx_top
//  /_/ /\ \_____/ /     
// ____/  \_______/      
//
// ***************************************************************************************
// Vesion  : 1.00
// Time    : Tue Aug  2 22:19:26 2022
// ***************************************************************************************

`define IP_UUID _tx
`define IP_NAME_CONCAT(a,b) a``b
`define IP_MODULE_NAME(name) `IP_NAME_CONCAT(name,`IP_UUID)

/*module efx_csi2_tx_top #(
    parameter HS_DATA_WIDTH = 16,
    parameter tINIT_NS = 10000,
    parameter tINIT_SKEWCAL_NS = 100000,
	parameter CLOCK_FREQ_MHZ = 100,
    parameter DPHY_CLOCK_MODE = "Continuous", //"Continuous", "Discontinuous"
    parameter NUM_DATA_LANE = 4,
    parameter PACK_TYPE = 4'b1111,
    parameter PIXEL_FIFO_DEPTH = 2048,  //set this to 2 power value of DEPTH = (MAX_HRES/8) x 2
    parameter ENABLE_VCX = 0,
	parameter FRAME_MODE = "GENERIC",    //1-ACCURATE, 0-GENERIC
    parameter ENABLE_SKEWCAL_INIT = 1,
    parameter ASYNC_STAGE = 2
)(
    input logic           reset_byte_HS_n,
    input logic           clk_byte_HS,
    input logic           reset_pixel_n,
    input logic           clk_pixel,
    input logic           reset_esc_n,
    input logic           clk_esc,
    
    //ppi interface
    output logic                       TxUlpsClk,
    output logic                       TxUlpsExitClk,
    input  logic                       TxUlpsActiveClkNot,
    output logic [NUM_DATA_LANE-1:0]   TxUlpsEsc,
    output logic [NUM_DATA_LANE-1:0]   TxUlpsExit,
    output logic [NUM_DATA_LANE-1:0]   TxRequestEsc,
    output logic [NUM_DATA_LANE-1:0]   TxSkewCalHS,
    input  logic [NUM_DATA_LANE-1:0]   TxStopStateD,
    input  logic                       TxStopStateC,
    input  logic [NUM_DATA_LANE-1:0]   TxUlpsActiveNot,
    input  logic [NUM_DATA_LANE-1:0]   TxReadyHS,
    output logic [NUM_DATA_LANE-1:0]   TxRequestHS,
    output logic                       TxRequestHSc,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS0,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS1,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS2,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS3,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS4,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS5,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS6,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS7,
    output logic [1:0]                 TxReqValidHS0,
    output logic [1:0]                 TxReqValidHS1,
    output logic [1:0]                 TxReqValidHS2,
    output logic [1:0]                 TxReqValidHS3,
    output logic [1:0]                 TxReqValidHS4,
    output logic [1:0]                 TxReqValidHS5,
    output logic [1:0]                 TxReqValidHS6,
    output logic [1:0]                 TxReqValidHS7,
    
    //AXI4-Lite Interface
    input  logic          axi_clk, 
    input  logic          axi_reset_n,
    input  logic   [5:0]  axi_awaddr,//Write Address. byte address.
    input  logic          axi_awvalid,//Write address valid.
    output logic          axi_awready,//Write address ready.
    input  logic   [31:0] axi_wdata,//Write data bus.
    input  logic          axi_wvalid,//Write valid.
    output logic          axi_wready,//Write ready.
                          
    output logic          axi_bvalid,//Write response valid.
    input  logic          axi_bready,//Response ready.      
    input  logic   [5:0]  axi_araddr,//Read address. byte address.
    input  logic          axi_arvalid,//Read address valid.
    output logic          axi_arready,//Read address ready.
    output logic   [31:0] axi_rdata,//Read data.
    output logic          axi_rvalid,//Read valid.
    input                 axi_rready,//Read ready.
    
    input logic           hsync_vc0,
    input logic           hsync_vc1,
    input logic           hsync_vc2,
    input logic           hsync_vc3,
    input logic           vsync_vc0,
    input logic           vsync_vc1,
    input logic           vsync_vc2,
    input logic           vsync_vc3,
    
    input logic           hsync_vc4,
    input logic           hsync_vc5,
    input logic           hsync_vc6,
    input logic           hsync_vc7,
    input logic           hsync_vc8,
    input logic           hsync_vc9,
    input logic           hsync_vc10,
    input logic           hsync_vc11,
    input logic           hsync_vc12,
    input logic           hsync_vc13,
    input logic           hsync_vc14,
    input logic           hsync_vc15,
    input logic           vsync_vc4,
    input logic           vsync_vc5,
    input logic           vsync_vc6,
    input logic           vsync_vc7,
    input logic           vsync_vc8,
    input logic           vsync_vc9,
    input logic           vsync_vc10,
    input logic           vsync_vc11,
    input logic           vsync_vc12,
    input logic           vsync_vc13,
    input logic           vsync_vc14,
    input logic           vsync_vc15,
    input logic [5:0]     datatype,   // data type of the Long Packet
    input logic [63:0]    pixel_data,
    input logic           pixel_data_valid,
    input logic [15:0]    haddr,   //16 bit total Horizontal number of pixels
    input logic [15:0]    line_num,
    input logic [15:0]    frame_num,	
    output logic          irq

);*/

`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Br7jmwnVpYaxd0AC1e16CFW6XhDkjFZfolVBd0LHHa/kpN7VVUJyIn/FqH+6DKNg
LewCWCQyLve1539J3WvRPmZ/ev3lsgHIGRk5U2I+zfjkkRnoxa6p60Q5mD5pJ9g8
Xeu8zUtmhlepM96EMz5eyeqVUuSLj/2VbBtSLMFTtbKvI6V5ZJpeqYH0vPS8XLVf
Tn2dPetIyBD8Y5Gk7qwt6Jqavus4rPm59AevAvhuXIc2SrYdEzw3tyK9p+8nqbTE
Wm/Jhm/X3MhoDn1gUQKol8mKg9SO5cCXXCyHFDJ2bXcfCVyyCSF/7UncY24duZ+V
MJqTYoOymPMOcy58LGxf5w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 944 )
`pragma protect data_block
2vlrkioOGhmplixP3NCJGxmGm+aPJWWME63wYF3SokcDRpk4+xgxdKlZblSRlyiD
sFGXJUMGipfVUszQTc6Al+9W5y8O/oCys3IyxbLhozEJgs54aS1Air/uAhMGThpN
yExeEnA+8qv5WNHEUadhpIV+uxmF1+PpzMd+33uo+MP04JhnwAvrZmtNmp/m7b4c
mV2ziTc/uKxLE0KAO8gqgUYlaVyemyqA+w5cg8hZ+XYtGaGIAdIBpx+FSsvhBGmR
uSU96YZ4rxlncirqb1wNvGZ+0k6j0K7vCswgvVzNs7cfIuUXfkzJ7LP9/eo8gnw3
2ZKbkt3PwVGGyRI8Cs0IKIr5+Q5ULXqZPzcKYuCP/AXp5h+KzN6Gxn1fwhFLroFw
r3JGzB2ZmlqFd1sCk7MZLhFdZuXUAlXlzpu2AmkObftolvL9I20DgLZy2+64N3ap
/p86d7Z9HQBJUfNuKOEoLa548hNhvhTUsN8hpRrfVxmbFIRVcVgBaYaSbfvxKIp5
Q9jLWd6i5zpqttuGrPJMKKH5WCQnnplZmybv63Hj1yJM1YiIihe4qV7Er2t21yiD
QmOfqJz5l1RbEZ8dMIN4RPgtOlera2eXpqFwqqBqFFeJPzwH9K2oZ3eWZHSrnPFq
pegfNKi2UtAqTucSwQ0dzVTW7O4u4WAOdkjDU1P68tGIUrnZ9OBtz9o7CG05yEIV
/b6apu3zXzk5plnUF0MxnH58rWlC2KjnTbe1rhECO0Lkw4DTddKP+ECUr949W/Qc
mkihtG2F2CaizjZE+a3jT7VeZTmYxOM1cBpbJfj6rDUWh7U0DVHRf3ZHaHwxAriL
wNId/274PuPNltrcTKgwlQf/y0qVkXfm7OF5yR94GRGCobSBjBiBVr7Jwd2/piOe
5Nf8bJZ3AkAW8GkJ+KplreTyvmSIfEUIWQlWhQvxddtFys7AbtF879hW6tFVj0sQ
brPPF9YoD9UAh57o9UCGpzFyvQdMZPm4NGpxOmdYFVM92yt0kpbelKJa5HLSV0JU
iMrVYkzHslWzl/lsJ0uwBOKbScIKyXGUQYVMACt8fDtQ/0jNvGVcHK/9/186bdlQ
zN6Ff9jLCALobR9t/vfAOHbVWqeSmQbP52VNExTwzfdkBi7YZkWXEzL4GYULBdNt
Ku1DK1fLYrlUZwakp5KWXon0m4naePWIrmEiH8k5MG0A1LfEMMcuUrjTw7qJT94f
Vflqxpoay05mfWCoorVcMFlKiHpDM1zz8YeW86i1KxA=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
gDJDNlP0yDDkgEURCzVzlCv7zzuvyyQ+UJLWEso+fi7q/kR8BrtEEpmmimoRsLnq
fQ9PmL73xTTNNc4MhEWDUJ9Y+6PllAvaxK06/hg3keYlCHX7EO9Yj6kCHUZecBYR
yH+8KeWm47TnVIMxQ3LHLnoEbqXMPHSI9En/ToZWTUeRQ8fLrbV1j6W5r7IZ+7y+
W+n2O2NeeKP5/0Icq5MbFHQMK7aD5E4LV+1HUjzz0ic/6Ge20xH2/KtuXNISQNYU
lESlYf+q7qA+P6yU9yeYK4YWoSz2p9B/YaT4iEC7MdVXXygurV38238IFxsapwl9
VYMoV11OcF1DU8O54BXI4Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 31312 )
`pragma protect data_block
lwYfU+pQtRGMRoCMW9+N8J1oIQrOPtU0aFWu/1F2IUTVYCxZhMkC8DqpNQbHngZL
aLzJJfXmsPlJ1uZUHF6aZarpfq+djYlUdav4/evILobXhVeJJOAa2W/rqTXC0ubt
d9P1rTOcoqXKEI7LgEzV5TpkP4ZafU4fMhV1dcRkCo5XA0sFyNtmx1Uwrfus3DrK
JfAyVInXqZp2F+1am8Ou3ma0SZ9CDJAimC+K32XE2MxSRpRnpU6USKeZ2nig+s3J
bWQpepnAjjoFT5Z14SwAdxQ0iT30HO/PGhCTnRwV9QMs4cvmtkoSDEhKKDbFWlVe
ZkSDCsbku8QmWf8dDm+sv8X0Bp0tGyHdNdfJnBaTnB/RZUDT2TVnvW8TDOp1Tx7T
bsnsMtAVwLf86cW9vYPJaoJXqM4qVDjtg2TTcodqNqppbcFVY0V8l58hWUgq3Q/s
duU6nN8y6GIuC8NT5FNBojhOLSIreW8gg+0fuQDAvJFMt4MaWmG/0UH2NGexB5Eh
SNikE6GdBxq3OcSzsFjHK5D858HK5o6bjk5ZaPantWRrwf3v9t7jcxYAYAZqo5Ab
lYAeMTw26l+xZ4xE//xO2s8JpoaoSx7CvYe8hqL3GLdWGR0zLbLLpG4vVyJNI5OG
6a5Y3swCckLg3jinaNKxAxCeFTIjAYouUBgQQ5sVt3s9e3O8i5JXYUgyfWrkqrB6
5yFPGd/ZdlDtd1uD1n265+EKsV+KTq+7AwxQDGbJdqDomhWgQboUxBIkUcxQQ65G
hKazXLO2GVo6/d/uCIl9E5oy5A/YA0GselvdCFBGR3RYuEpqFzIa5neePGPRNyxK
SltM4h+nJyuk+rA4ugiKLpxyQ7dNOsEK5me1Gt5Kblktlu5K7anaqUb1/I03Ji3Q
OXG6ClL+HN/FjkqLri2uqd/o3zoHHgo3aRe8LmUTZD4KmAonOp0flT/nEq2X3d0U
vyrkempfh9vAfimvv01AD183Sm/+XzUq0Sc0SVU/pm4365nlzZsGUKPrl0F2yNwc
CvKT5z5Bt3oyWpzSa6B8Jz4REcg2fI9TuFUGYDz+2rih/VQ8eHeLjb4f3NkZqDbr
Y9if9QnYBs3qV5loKc6vzfUzl1U83V2yHeT+dFP3xdNzgLnUQ9HZkObbtCpzCZTz
gU463qRouIE5IfDarBCXucLgAQR+HpHWEBeRPlVG+IxXcP3bd1iXLZaetf2qMpli
7ia/h4NN0bKZdu2RjFzAqA63ZeOTl30rkEH8JmaV3Jv0Ftj82V+z0eNqPWayW0wE
vFXeDvNBL3SIeUNuVr+N7pKJhQ4mMgRSDmr1BC+a543wyGC3ueUPqi824xTumZVI
egMws2YCocQG/fxKzIAAIee9btoZ6MqPNHwIQw45TPAsz3Afl0yx8Av+RpDxssnK
softvXX5u/jMRUgAy/2IKZ2jFy6MZEqyKhdq/s+Y4NWWgJOAQ7Tl+n7pWpIiM5Kp
LPaGSbsrLVit7LLOWK3f3tNWbVkfJ0ZjVRt585J6PHIhakWmTXt4AVj3+Ta2tc7r
m0YiEh0pI6YKFr3WXrAqQy4TmZeF9fMpjgu+Xwh28lM7QKBaUuC478TRfY4fj3z6
xErPj1NbfC0sDtAnrSkJlrKHJXPwB/A19HhYldfqINENlG7dcBCh2GBfM4+SYWD7
1PEyu8xGVIBfA7jHBbQnP/zqJ0362PNyqbMxxOuS26WVHbhNhnnVxSfHhRitpyRj
IUXuuKAW2arsc4Nbbkoa+8OTX4JPJJenO/unre7kOik7w6/PPfjTWE7xMb3wu7ex
/sbDwJmFzSa5etmmPQA8ulAn0Z8oJRTnfiJKB+jYQr4CHe1Op5s5T+xE/wUczz9D
o2NwVyxCE3UtfpMtu4Wwxq+og960fefA/Lxawre71YAFdI1ZVqPHhniu2zsldZZx
BnUbREEumjJL7iZLZch6Zt7KVwUll4fiOqYC4ygSDdDqWQ5SJeavSClAC+GqWx9d
FqJVMnFF7dlBIVRY6LsJZlfkTePXgWw7qeJfikEnul38xxML15tYA1XTh0r8JfTG
VRxt4wvcXQPpG5PMcACTFHC5x0jskaq8EmdteJBjhGBPvMlv1O5dM2BC0GXbqdGs
pQJe7MbqIQzsNfsMkUQRCQe6JFQYjQ/LurOvP1gofHYECktP7WKWs+ENdwbFbGdf
PxZOA4A7GjmrmFlrgigxEbmtfARYFKm/qQJEgVX1WsZehvBd3HWNQDzBeUJFe5cs
gnJpWPZETkzlLUc8oFoa4sfQLerwQ/NH5thkY5tW06YDDcKoT3H+rwy9s7szcjPg
cVQtQsE4NhHnsB6K2CrVRok+NYRfUuM5e++1gu2zB/RwSOm3oeJyfZ6NYY2/jf+j
y+2P38FsbNMCKjOw+TX5iktz5CsEpqLfMFAtE6azX1H5H2WEJv2k7pCsCeqVMQSP
xCOkTeUzZ74nHWF5735KsyJTbuDWHkrI/GeBzKOy25CpxOeCLxP+DJs038pt1Pjf
ufRklYI1OQSjmk4zy7AVbeOy5xL7byDbWl43XUnMMkDglMGxNTV0nbiwNioXQI2G
cZ0bGAooGqWykfaWtcXq35Tw+iOmI3bgLMX43AY9P8E0FEZN41XAxdRrWcRc2aeO
lvUPEsoXavEsUf1i5B4taZrnHGYKnL9I+DIeoe76FM9jzdqFz6+JuyC0arw6O1hO
+UbZ5O+wEj09SqalXshwPvNj2Z65eR5cfpwdeDmjJ4owGHR0HkaaCjaDOXMHxJtE
6GCfIUAryBcgHhfVdFnWpIdXBkNSF5VYIsyMm/uDYEpBwFuVSWdnpZCL9rUerkpm
YXom2vu1Qtnyy2Kh6sMnfmZPCMkigZW9ySEa5aedS81Uo1/r/SwcmH9jew89TFJL
LtaHyjgsyAsu209KTTDJAo/oOcjvd/S4oeHpp6QuMW7es3Jwsbz4aTtC4QznYYcd
h9k6lmUeBSpokFc+lAs+IjcsF8yNsMimfEB3sMSDsxf5EGBkREzDuy5Ez0fNYO33
dpJ1U2FvHW3LWMxHfSgA7niPi/Rpsc2VUKx2M7iVre0PWJJL4lCOWlJT3OfDhpeq
TXuN79b8E85DvxIcCGHwxZJXwXMqrcQJkBAFHdoplX9HkhC+VCdEv12a1fmNaQnu
cZuVzqxD0McihMRKRQDWCRkP2dste0924VO9JlDsI041HpI0W8aMz5yA7ltNQ4vH
14vmshL90bK3ftRdbN6N7Z924owngJBxAfUk2j74mvdtyoxur8UBBevauh/SWS/a
NdAD8zhr9IhfHX+AwdL/fCOahlCoquqYQ3pCo5AjtCeZslDIwrQlJnERKgPlBHEg
A0x8XWNuyKvauXAk+m/TNN+T0hoiId5bN9BtZWLWt/5u1k35M1Rs24OQOC8KXZI+
Nmns4WtBEGvJ0hGs/xZmzKMCvSw8CIoDpPMSDjPIQ+/q+8/pncXxIB5n+Pjk++Yo
vBnvVUADnRhHSs9qG1DNFXI2R8g8beskUNqiB0q61NF7PWOoWxbaofew9CEZj9pq
E/9BKYuhe2PIlqgmZWDvFI5jLCqZEXqV+SZH42uvARchgSfPk1n/9p5IZagawulf
+rq18+PBKqDTDgv4zrmeunFiRwJBszXdZc/mUsi0LuvLajFtE3jXs9SZtl0cPvqk
e+LNRk2xweLzBdfWIhkwRhgMIcpmW0slDH8nV43UjLEom6cw3SIj3vZXjK+NbBdD
XB1GtLX842aJObwp57ih/zFXzajWSDJXiWqTJl2xWj0DkUdG6pM9DxePwWeLfEya
CHFyATxwVlA+QykmSxxet8IiBp+iFi09GP5co73eJR7c2f+a2YrhVGirtk4LTq52
D8GaIBtlfNOnwBMZVxiLvSOwfs1yyIYfDaSB6t6lk4VvDpjtbd1YFPXd0PZR6nPA
IWZYN5rcKDcDPjUn/GgFQxHLFCH3DqgekWuwlHXhgGUIS5mplH4tli0rsWhHiFFT
StQAl7MWdtircj3YxsuVjgHXEVSSAfdRSef4agbKi8WlRx/0AhLf3Y/fi1mldn85
Z8dHmwAjqqt0D1GKks+bU4XBykIvjpKKHtkPokTZ6Aca9ePF9Iffw7T6eAM614pq
RqAER6fFrgZID6BgoT3szgCPWSISneQxlERFdCRK0VaoVCZPxMkkg5XBCv2LZpD2
ELmprjPUeeMVtuYDxO5WOfMeDBrG8z1zyceAdePEuFSIgU8bDNRsY5rvkxmUYTZk
9sDI/m7aIi963tamE2fKxbIVxEeB5Obt1diTEb6ctzskfkkT+Sn5HAxXLFewfZLG
jGTJckwBCj59BMEGC5jYnxYdT70+jiVqnR0LEf4y/joBJ9/lElDSVMrIvCFqcbpz
PH8TjydOUu5lVPJL24vF1s/kKyRGcgPg0VPfv5qVUTHjss25P0fxkduHcPeRy8WL
KHUUlJCQtQDoIKMudKTovDGBpCGbNQF3HzFMMLOl6ekgWib2lHuueFQaCYBgtVxQ
acFcr8DxtQgeE/VQ4t2UCwccbVEsMO+/WPqRKDeq8HrFhmEkYRu1KX5pl97o3krs
U1I/21jfNllQCP5XO2h71YSzWtS49QlUB8c9kyo0jH0um9O34sqGx6zmwk/9Yja4
AiHmvjWDlpHVLy8xsc/e1Y8AkC3JjQAcipvRi17EMv5LPgCNBSrzJ1ahYlycWVhM
aZvMst4RueSlgtr7RhxMGlRfCKR0bV60BoiTzbApjCfOrhKWAGtNRI3jT+WnxUre
phDegBuwUVPkNwRPVfvAXVqbNbEDv1uaRMarOx/lL6XtrwhQQXQGi2WcPT1QtvK8
SeNkvRi+mbFymuW3xnEoKbZV30u+nIs1EcxXiYBm/0IBc4XJBeEnBnMbBBqr1hgX
bgKuzSOxagKbGw561MGkd5KD1LoRlrJ00TcWE6BFhiiLtxVVzBq8BRzjwBbOPYPn
6yo0RDP5g7Ygd+K/8YA2zVonoPogsWrSeQkLehP7SmqHvkzv/3fhKdZFAGQ7/zDL
/FA8YVvbwnzLHn6a4wR7Qe4yiywrtX1pneQA8tZ2lqo7Svv0wPKBQolXq5suhReW
CYeIb22O4L/a+HLRckVFNgOx6wmNM5K3uDKp56Mhx+X+HledtZgkitd4/Wte29nY
h6oyfIltSvz3LuL72/EZhqjDsUXfiw035+tyt7o3NdwpFHnVa5Wy7fOehJSn01xo
vHOA/uk3WWeo8M2OcMAciS/cYumhKIf2By2fRUdco4DpACadXxF1nvdw1iw1Ee71
+S3AI3gKk3WZH3lABMcLrUbixsO2JexDOSlUV1yhjP22Lo8TaHHRrP+mypCpMjHE
u7NMXV0rr/goDdl6zwdrS57jCqWxxrDsiwt+74w9ogSGDU+JkGTLVpWAW4BIZCdr
JF5OUPDTemkqaYra0SpAU8tI3dJM7j+kMOsZd55Mvd7D36m6GG7NAs0nlwdxEoK+
22ErkpOA2EWgbSbLfx89vJEqVMxAaGWpblck2mjpu49fKwM/0C7VL4b+fANgzkXw
SyrPE9ymuUy4FEJElGisa3w4MLRAdP80yqTjKXdsHT1txCE6iaCj+SnX9t2UWrtP
WBePGuev9i67IZOvkj6AKNTHfdLD7/PWKHcky+kNdambTH9Ff88OdJBLoZjdk9vw
R88OP7zJ9lMfw9O49z3m+YEYY/ZzzlQLGxHgzfYB9xdcxBZSTcHX+8hIJnDeJiIU
5qjfqmEFdmSJ13IIx+YYFmwpDfRFHqlUavpYvirVuxe9wlyBV7oGTeuG6N4BYI0f
QDV/GGggMdHmOG3iM/BETTp5AHUiAsYXiqdFrmf1vDUGyz1saMJp2/+UhcqqrDhk
xm+KcMW3V6DMbgrVHwJZp6Vf/i2491HKptsY5ocSRi+gPSuKKEcg7mzfWGIlpe/+
pcnMWBDqa2FZu7wU639T4TKrlzrIblmt8O0CFyiKFGcM4RZH0DI/wfeiLwp+6gv3
VjanNsU9oW6GVXT2yWiAnW12kWiazq/0Eh6hSHJ3oDKAK/2st2KKzoyyJDSHWDO/
/644Z5VNzDOuj3AgZiGynGvBh6ALs2gkn3Nj1I0wNUZntKYP/0Ikmx7HheGubMzj
pAozYnJRbaPcrXmeiTZu60nw+08dqoZC7/i9sXhorxRMKX6kAw1FSL2Mlna+S9Ag
UHz80K6dAQ66TbIp35nroYk4c8dcW/e4a0riB0QK8apvG1lNR4LKWh+lRrtqy/eA
6XfJqgH39GDRyLYLq7tkub3nLx+IF8AQ8ndyXeZlzlJLMDHjxpi1JPdGwX5eSjdn
FDYO2hRHvLn+oR93WVQPul+/+lv4U4Va1zj8QoiHAxtgiDdcQSceMPqizR5FGlNa
vT7wCzIecspKb4u/4Gz3g8JmiQN53x1c31GtLX3IAqXbWhAjrTjhhL1x9hi6yw36
KY5h9SOzDK2XOj+lw79at/TmtgEcWkMWxy9DCImavKqAHQr/c7nXpSGxB7w7JMXN
VprR/XxKVsen984zoZliVW2T7EoPVpK9VEH79T09Q0yAehAHUJdbxTtmb0vDV8sW
1wSXIN7BZRydRPI21rVJ8VwyS72+2lbgWuiNtyrkqCYtQFsQ3/KNEUYfubZfg9/+
PUuh+hFDBO93aEnzHvWwnjE2zD6/dCyhbXRg7iAbbJssm2A2gSIqapuETadMX2Ac
mFmjKYj/ierugdjsa1BXetC3aCnGlWgc+JC/tF5HAHRYhibQwLCaj2LhlqYuX4UM
O7rUhB8XVsAJFVCdPagEzFmAg+wK3Y+zZh9HoJAe6cydd9LJCjUuXRKQ+hxG3PZ2
FvLNpl4mH7VyTI1avutYAuIaJ5PEfhsgsIiH3DwBAyBpZ9joHx0Goucj0iKOLrxg
sNxRd0Km68ubaHi0MZhC4pBw0s11nJj0PitwfA73UVpyEn/RLdUor6i5p9C/Scqo
C7rLK1vXG9g8XryhuPdLenPih+ytWdY5eO13JC5Lz5hCdbCAkdUAVp+6S43y/my9
k1T4/qsagQQdDNH36NOZVanwx6TIrkhxXO0pxP3TRn5cPankKRajoRnEjqHjtDyw
Q5KKNdg3ufTOlue55svQE0O0dA0T7eH3N4kkBQT5z9d3wKBaNrBI/tnnQTPR8fK4
bah4l7n8wwSwP5UoRv6gedp1jCtLUWzvwgsTPsu1QR1l7OniWFTdz/bvS99WdCoM
0zYu4ekGWinQw9pCJSwXrk5PUztme5n7GcUy29x5Q0Rz9L80ydoKIUkLgbvHWmaa
OFMtuppV7ZB6DPxlNLAM0x87Bnk0Wllza9Ul1KmjF3SAAZXgmAB2trsl72C72+Iz
GX5bDwAkmAvGdGlp04Tqcf/S0IKlVJO9oqwVjDE3lhXp+EqFty5KS3YuAyIYTDGO
ptOd2dlRLi9kDA55kLttKwjPdyyFDE93ZVQXEdoLWzGDdpwbgdlvtn4oaR2getKY
sjscs0c97vZTSiiJFb5KhMmId/AFb9NKd1Gn+bByD7qpCwz5+dWDgGtOVfXZkHcy
8HgbS0+cZpCBLMIxgSiRA+aFirZzVGpOwrHYedw3xQ7Jnj3nSxghmPdA3+ICvPL3
PY6G6KTOusEBUfb2f7jP7l4CA8rOE9l15uqT4ewfIvkg1f4g2BIlwLlDp/3Km2Lm
xffB87NaHZW92gD3IUU3RAdYIXo1sMUz8oQIGwPHMeYjzBCkcZFxgOWwJ9KVLVkq
ompOVwzcA0yn4CbQd/5QG6ZYvYdEBZlL1djuirgaZ4JMDGEuvDcLe51Ob5hJI2D9
CUEwr/2enEsyweOH5DmqfvXNOadWFTtM2XmPS9Jk1JBj5UpaPYfNIGIv5vEfpl94
aQUj66e44X78urBgYSP7dGfiDWkzAugf9TaW889aFyStJwPJxvLJnjsR+8GsTvLk
i5t/zVsKe5rvIcfnCI7F+F8/qU/dvu6oP8yANzdGT1dtGR4HEgjBESRHd0fnBFWB
X8P/lg5zdsf7spmMi0uhu54u8kQk+3YXQo4xY9ieCjUpGIIew/r3dfwm4ZKryYg1
LCpFzXF80cDqaWg6+BDTk+ywta2z/ZIR3QQ59sXNL2h9s+4BS/5e9uxhfS2ewoLJ
IZNmhV36Me+me65hMsyxj6Ee1RlR9PDMwrEfN4uVeiVMeef6R8L2BuxL2F1HmluD
C8gXAVL9XQ/F6qoH7UQ+7L4JaRkptW2UIj9s3uXgZ7U8DH7NIrub0WGR/J8hteJw
1LEltqBw9jTWnw9jgcY03tL4+0/F94LkSa7wLD69GDz6m/GqB4H36f2oU3JuW6Ds
zygtvTZEgZqXUAyFharGQ6/Hm3W1lo3Q186ZQuRuICfMwbXkRASoWK+gDwqPtdPB
LElL9nL11lOie7bPlIihSROUJgZDrtYqCyvIM1a1s8D4JexMEg4c/g3L7/K5PKKz
alOsP3t5I6SP7/D3fkgRm++iJxO72xlW1QMmY754R9lv4SAXWh+0eA8dN9S1Yyr0
D1+ChpPKn4gutDeiWf62i87iMwcG0qBze7Bk8MKPR5xMFO0w2dHaU4u81KpLo++6
OYXMaP9mmBwfzLA/4sbZtk1M5hzdKAObXLDHcHksZ2BOoCt7aMDTThssOCpShTne
qibDI1fhv2xfoSRpAEjRYlgEpJBkUEZ5DqckdOzoBgKqRlUWJM7UStWh4zKuAgVE
zBNTl7hjV36iPRVwDOJRHda96FhB8bG1lpnRwTpOAXcxjAB6UWac+ZFkkzgHDwmq
GgSN2eXhGBkOrdqkRuO1Fny8mKs4jyyYWC6tOIJHXZnMvRZbniaAGcEGXFvKl6FP
kdS3cYfejxEsplUjuzEV2eDeEe+BUYS3eumpgVWm+NeYh1XSnIlHWM9atVdyQR9O
JymkvO8WW85aEAfuFggOv1N6nEk2xZZ05I0mx+KjLfTwb7L3DVRa2MocZl3nYkzE
m9UPMh7NHTTjRyOYBvRKvrdkBRkxcnFrkUvdyoyUd1uuq5BiqGhJKCYBl5rCTt5C
4YKaou3y4P3U0zNfHXdim3UVgOCeSRxrfOJieyodMP0ffy215448g5OL5h9zIu32
zMIch4Xac5j6uX0+Se0BYgS+iH08vi33PAX7SroCe3ZoAeC9jFC5xY1SktQgaOtE
kKSGYQgoubYgeHTTD7Fj+QoR1zNNXChpGkz1NWaAO/Aofe9AAExQ3yVT7RQ9VsqQ
VY5xnqz8qM5q/pwsp28sY17kTDBVKrh7P1EsHHPj3Y22rFr5XSenKrzSfnOqIcsv
vbX1HJ+h0Uvwvvk2x5vpZIM0jtC5X8/TI1lSTaoeb04+TyD+F6Q4+9/cCmwo9gp5
o1AIfPNgF1jsrk4WysYPfoD5MceCUd2JHyjs4oCJed1KMw8RGrbzyIbtbwSdo3yR
zgOnYe506GONKMqO44mwidBHHLc53t6kWFSsj01Oh39g35dnme26vyttdvSzd/lF
gl38RM4KTZkrV8R5D2951Pe01oiD7mC9JowBq9UcjWuYAh0oMBy6RqV6c7mh9GV1
6l5Ts9gdkNkznPtTo7bn1bUmnte/ez8wBfEBYeISG30jlnO2MNFZub9ebTZOuO4R
pEsPxd+ZyID0eVkboyXRRQ2XHe1NW46Mjbm9mazYqf8YYI02JP9gfKCgxfqGAiqQ
idiTLTGl+iGcW9mTricpVFSSjoYMnHOUs7WZ25KT9mAvEoofoJlm66cajR6aqbpl
PSvKSaOEHndS/OjDU3CvOcsBwukqZnQK7nPsCWuvwTWFb3bPb2uW1niLihJKFipt
RN10KY5HYUz3rM6UffJXy5c9gKU8BCkAb/SJcfIpuXIZ7X1s0/nwLCojSv0MIwwi
xc23EZ95cKJ8sZsdHIr2Gw2q5eUtW20cfEpcB09gn420f+sVFTXvj861jxTiZaid
Dq5gCj5rwhsnqPrSpXNebDOW/nqnGcBfhYu2X3rnLmT+K0jwykgfTAruA0QhLfZH
4lCmc3FVQa7tgyIcEXjQ+C1oNPoY6j4qffq4eiQOPXW6NIOVMRbhTz7P6dPpoUSc
eR54A7XXRvacgTfCSbyaZNg8eBJY+4434LiMhbQBDo4+e3uGQUQVoD9Kdz7Aqbmv
wZLPFMofGb/UjLbXYuRrr5N0KHJ/s6hCVj2n4dlO8AZcycjKDNkKyUQpmB8YwV0n
BIVF7T3alU6+rAsOf7KXGxVU34dPelvHMcZioh+Xo/8Euj/kf7SP7Hsv89+TAEY2
lE4Qk8dW0fUqPlICdUKzPqntAzkNmFnRVHq3NadNuC8B/ipTZvjyRY6wEJr27a19
hi6H7H4O9CEnU+AGs566FJ3IDfuQi9jcuW7Y/4Zbq9a4fr2iB21LNQGzx73iveTj
6bSbSQP9PMPK5Ki8XQQFhOQ3oGCDebco452ZNTxOaDogljMDEzsy3HoaWtD35qIG
IqOOO6lqjwiftRevNmTghp3u/mTJ3n98a4jyfKID3z94SKzXRGjNe+1RH2GxSZL4
6mtBRLBKcBpnh4+YH9VSXlG1xRdqHnvRmfZMhObsl8ll1sCYey/oxzrl/1QOkDWW
52ZdM+v2lED1OSbi/itMEaP+R7yiNblLRFeVGUuEWoMrnPTZGRSO6/a9b5USD7sp
RHmq5MFb12WUvB4bbLKcuS78PcL/I3UD3u4KHMjtpJAcj8e2Rz4bg2Xf9tZfsWZm
lSCH9h0aYd8kOeozKPvbeA6QlIjfsuSRM+oVeYY7Yqu0iZRq8ZFIj2WkAx/Uq+Bg
1nZ0vbeq+Up30xaNBgngQC9ayDks6np/cERTvPreQx1IqM1+yOnctrwNH9+KTzol
mtv4gICDm6S6h9oB+z9AD4mSqjb/Onj4AREMzfcK0WOh+U/cp8BIhrKwuLsRfEjf
FQnTAp52zXItkXN894OFhEyinRajjdmTZCy4lVoZC6YadDSeWdfNsWuMrsY3k9BT
HkgpkiEk9arvNJPWOitfvCYtOltVIC7M1Ae38uRMkirobARRvgv6yrPR5vHfxqu0
T00zM5j+d6Vq/x8XWS90jV0gl6y0mseTayPOQgMWodIerVAbGR8ya36dzKc7dxAJ
M76kXYQXQRqpUkpt4Mqn+/wCkrwMv+Ph4pDMeDj9/K6R4p2+RMO4ceZCZFjaT7br
bMiCIhibk1ax5bjW7hChbK84qYhFUCgFqt4Hz5IdZIAKf1wYi+AkF7b7EsAwfoJP
82ynea7sJVg0Qpql9Y9cI2XfFTbalC8b7vSI5z+E0nrpIZAuoerqRXqGcq+jJ0Om
ugEgd//tylOS5exGuZ5w2RtT3bWdj/KegTAUJ9+fvCQN/zclQZOB1FWNgnbV3rq4
KqYMKcPmuDsEuXGtE5pBfYYCfQKRZEJR+JRzWGGDpyUc3Np0sLlSPcWjDQBfDrkj
XOtXxfueBrTNNA7KRwmAkQW1oxpftLpLfHFUhv3OmPBZ6n6rDmNL8YZ4sl8tUzn/
FxF1q4/PZ7cKjYu+/8i7LNjySKOdTiTYJseSH6vpMOnJH1+KKYFg1hdi6DZBD0u5
26ncSw5tD7Hj3ioiJYkPvLkpJ7BRVJjWyfl6GVPKh1TN5NeWGX7wDfNX/iwDLjPs
R1kcp9nI3ZrSMJd12xEaAL1N43C/btxjSmBMqyDF7ERlFaNiJlioTwd1yhyLVyoJ
iLSS36+krWvHyICVntHJv8EaSJhe4Q10rZrRuC+uN/H4lFbmqHnqFK0BlBDeRMy6
h0R5AMN/tAcAPEZ6qLyr3doq2fU9pjOjrDl3eEt5sXp70yHnaHpkyRV52gVhzSL5
dxRPJ+w0EFrajtAEIpWIcwG25syx2kXT0GrTWBPFq9jzqEVKB5IiN3yexf3FL9dU
x0shMYaVBZTG1NIS9tMGWuBnK9ahu01ciYL4pfxv9C8e58nQiyJlT9qdZ0vAyw85
bcLTCHQU137pfGfrJkrjm9Rva1djkBINtmwIeV9FJvR3OgazMXk8gTU8/PZEg7Jn
nNAgzae6ycEewX+OAOIhNgGftUOVSYY+NFehh5v7O6/or6AB0lt8Mi+vQ3nSpdWp
o2ngpkosd+/EF2LUZjycB34BgAvOsBRRmD+MOniBMvcITey4w/wcgnnhqlwjgoUb
hTbyIph7LZwxfOpZnKltmM2BK0Ka2kQgJiNOpNRJolHZEPIfKR8a4xz7lgkqevRi
ojWvtsfIutd4/wcNC0kf3tHa90HHjII1Cm+bi/FEo0A7JX4/VV7UMNL8NCnb2gSF
ISN/o4vlsvLgFZ4iD/uQ7jXm+1vMwhcxQpagOxxdNcbhzTKFElBsVZin8K1oUzvQ
5XbQvBLRZrh3eU1g+2S0EiEdXiraXBN33VZFZXrmFyA/JfC5zd38a01AS3Qy1v/w
Frl2EsLxTqDkFOBIpfPFNFIH1mxbvJsm1mH99jrwyrzuTBf5g9eV5Tb0FKTsn26A
Wtox1WDOrijRVaBXppPPNXcRDChmiEk6S2Z66J8D7TX4jgx2d+cvcEvZdNvvKkgH
LxGzW68nFjz0tGOgLMz86ZTWHiLsE96VCs3WPbZO0MtviGu7aGobpu+evUOsPtLa
l5Qsnk22CU3Yl+r2WxuR0DafsBlzrOnH8F8cx9JeEtHlPRIaSVKJt01fuBvZArBH
2vd3urs7gXB/mPIRA/m3AR2zeqe+6q1SYIhwXMRtIFxYxTlIE/EOLPFg3XP0r9bh
6FqQBUpuISDcSHRhUp0snK7xsJgsnRie8R+xyPoEjzR8nk4H2iUII18tBbAFAkE+
mizhIITaAi568PZLSxwJbPSKYc3y7tfYTWJcp676VcYFMK/mMsvfQQ9w08SXHdkl
1FzbAicGlpNxwAGqKgU+fk7iipsaYyITN+bHI3mO8kMr1r16GGVf5KEP+Xoks22U
3rIexcktgqAVW7nhmvoivMV0beJYz/WcJ/UoaO+SxANXjLThx/wdyWE3zD+OEgBc
FAZwaSQV3FidsW196xNW+Lhxu071bmmcvHcRh920zpNpHQBjaNydmSyaVWE6OXiK
Rdk6Z8vmETO3vCcWDFl5eEiZBEo7HBNbFMkvytCYX3ByU6a4VkliLg/J8L73E8ce
fKV14LuNx2uuT4sFCy/Id+/N+pb26RaggCZjQ/VNBbF5t1iyt7ZPGCyPreiDeEKS
3Ls9MZUJYRbrZmNcMUEsTOHTjYyQw8ihxFmrmoRzakVH1+FuwDdtRmzPZnu5YCU6
aMA4vw5d7hh/0V9V87xm+UjDUb1Xgb9UOHp6vFP/VjheJ05yQ/WDzFPnJDRgDLft
Ht0RUKuxln26MKW9Xz8NLN8yY3YZdvIzyX9rjNx3C8ajwxJx+tigPDoPx8tBeQ8h
yDRz9/e4Fv8SqQai43FWszBptg0+B++kVmg7UDmQ42+HgmD7J99ioLw+z7jhN7YD
uHU+16B1ZQ0fbXc8s5jplUuA+a/jzK21ot+JZOsCeOKktX62lkgfSHxme5l2U7GV
qs7kyhGfhkV4nst06SyTILxrT99LGadZi0xTAW9az4KDy+s9pzAsDQnj4tyK6F2/
IX/GvCPhA6zLPFUrp6O0xNhilE6XLcxbT135k1qWL8cXXVnE4CS4T+yG7DkVX7pO
6jXce6XFKB8c4DulkwuiRjXfZRlzc8EgEwyTKxCBiBMqgI7wUdjGsTRhcqa3DnIe
kw6ZPYK7tD3lkxjPu2udrH9h69ZujMEMA8Q1t/ACxb4dkeURiuFKmh4H5Haci4Dl
ge38TgnbWjQ/wQ7paD0GUKEj3RnUixa1jtmiAl8Jwr0RQnicnlX2YNQ5X3q00gPi
bk/FJsVo6ymK4rfVgPb8TwzQix0Ki4OMr8uKi5k/TJa+8Pp/bwibo9i+sPIL+Q8E
h2My47BoJY2oads2ZL6LDEvMP6TDBL+Vhe1exLOTaPq68NQ5CRNRsK1boNEQqYRG
cSYRbqutNMdaNS/yL0T4solMg+V4d2pPBERPhPv33SwlxGvgVwYoiXczyqr7W842
9iIz78DL6alMkTqacPaYogSmuDQuu8wR4q1dLfXcG5xyg0JSSwXD+YIiEJyvuN4+
NvZRHio3fk6dR+GYvobQWVFk8pPPnhM/bF/WTkvDbO62eTJlcJ4swlRL9gm7twVZ
ZKtvxH0maTRGkmKBGmK6yF63Uw/qnAYsPsKT90HdX731QSWvO70hXR6R2OyTzCoC
uyacl+1Cftbp38wm91ywWLaBwetApoVLa5BL6BT0Qkk0KydaGVtXyxyKaK9lhhlO
NbGK86XWYRpm9Ne4uIMuKwPnmL38VpYgtMO6uhAay46zW0vZt3VVid2O9nQrOLJb
FXmdywEL81velI7w9O1M2dq01QE+Td4qTbliRESpptxPJiPkjk0hs9DKSZgkkeUq
KNaUj9WK21pkIBylYymRlgjmRKkxO6QNP5DIxHzoMZUsnUI8Ae95X4IbzuxRHH9f
EEsuuSSDljvpG2xHgzRoSoj8hlZHxCE/yO1yvqctL6herlQuQulESWySvo1AittU
7G8YJjvmhn49QbGylb+b7OFDhui/fAKoON4y5ijjPXw4nOWjq+aCkBUputHPrkas
DzoDILF2ItP4dUmeMz4j5KZLVVgtL2PxHxQguAt0ZPs1AndRkaCsW7/yuPeK476m
OqWN0jtqnBFhKMZZ+CJHaIpT7Cf791gb84zCG1fIEcGOUVAT12W1aDhQgEXPUOvB
5kyen75/gi3R173K5JHGxAf0KD4gXIrR5w5KoU2p0WRj3kcQFYC1pPpnEC3hICtS
cQMdYfnikU30bECCWfbiEs0TGMZuv3ho+FuAOFD7Hfb/eHduJ8pFxOyHqH0thOkT
uCco/w7jj77q97HyaqE4JZJMCgmGAARgj1k7aK6JFQJpDpvxtRlfn4fcNK3TTbB8
c4NCzGVcMCQ8qNkQo9rm7HQdfvwtWQqCGedqK5u9kxyLMGFQhEM4cF7yAOgCUlLh
qrULCrH+bgMY6YufZgT+4T/ABOOPsW9leLM3vKBP0uZM3i2J8+gZYk4F91ArSL2H
4s4W45R8U5anbqOBMncXF60+euwIxZcYaU8Wam9BrmI7y5V1NPo5njkBcEQ9e1NT
v+O7FquRpTqBk3ni/9kWk9yNfYX+CJ3iqt0kYhjUbJ+2ikTzUtFmtIt3VjOAeGFP
wm4MPuM5+6CD97PQ9okVOBbpm9dGU69wzO80/AE/lJdTGqWtD/AZB0sDtRDCEPFF
8e/JfV0B7pnzUx9Pkdc3CJRR2A4WdlJxsOWHqfo1n9LxohQOUUbW4sQxu6opvD4w
eYqQfBh0BdmNLM2EHI7zNVU01XNNrc1Gm6ZWaW0LSuDwHbQgyLqg4c/d1cFKrby3
xam3hHdAjVnj6x3OyOSHhdetcnvlHPXd6IMIbQG9J6QD+Gqe+jQ0aHer5gU3UMOq
kWZzKEED+9j7CUEMcgbO0/zIUv5AluX5hs1AhnJNtwuWD45K2MxyIGJMcpqurTyI
UcFlHBeWBS+y1mkvfOb8FhWx5zz/jf+09Zag90DtkfIw8ouPRVzyBSk46g9XCguH
9jSk04+sFdrN/11mxHwe1zg8BZgn5t+dVvC1FHwKNd+bl/SaleGO8XiEpSaNLZv1
aXZ+qnDCX9HLZQxftQ4o+d6cnkxzcCOEHQxbn7peab5z2bymh/8eMPq0Qx83WDB2
w96doLP6Ma/YwNl9cfIbH6fD9dozEmGh18L1oQ059Ch/f8K0mszJ8U291R56uGBm
7GXpl/TYiDA9EyLlC8gOp8ZGJJ2ifxwzU6aIQeHse79jUZLOf1WfaXDLDwZtOlNy
IIskIaIaCaKqsLM6Ol47M4+y1hvucCfSnBQWrT8yq92z/Re8GIBSkz2Na3YW9lXR
yRkkdzpekS+qbzZmPaVevwHbaLDHJdPvMYYBgN9Zr7AvbABdXE19o9iMEtCemtQc
RSbQbX6PxMu5rgIeYy7BNJKo4uI/QGulyM4M/LZAgX7AfmBgQWK8fhq7bVRSC95M
DODERfucYzbptU4J0lfTuovejzEpHRW+hB8zYOGeUDZkh4y9QrmZSVdcUvv4l3/c
7x/CSByxb8bRZ5ZUL8m+UeKSuWw/k28nyNVpouuDtSECNqHRXEAgtxSYPr3n9WYz
+gqHkQrAoL4i2mPlgypIcJXmfzjnWF4Iqpb8iMdwvFs0yteoOPRKYjn+9202C802
PTRqRovTNKQI+61Xa8KwAjqPpySTq3BrRxmwD9CsGlnLTfdNwCRR+X9531HA8Xfc
jxy5gpHDg4Bpnq6hTPtp2FZXrzVmcEYeoD1v8QJLGK+Gv7y1JgK8gM7pWPktGLMh
F7011QXibV2X1vOnGt8Eu2fIZf3Zqo8cUR50DdX963Ni86s/opr/NOQe7JGlKL+8
hJE2XJRB+6mSEBRMIPrPdp0G7S+chlJNG6hkPvAYQ4esvAw0g4VTWtJ0sGSjouCv
T2XNSLZ52g3uih3ZFVYxJHub8IDaLyPJP1o9e2FaD+CFQCVO4vehH6PZSFgOFdbC
byHD9OsoO5OtQTpqwpD4QeTe7R43Ceeb9lOaiWOw91Z67ZQQvqVMbDn/WLftJtRE
05mopwUBHL6FUR60SEkQ9eTtjhfHcSBW7E+DlJMgvicph9k5+JfZjusDlZEGiqAX
XG14Ess+1PpJleDhCL+FIpaoXclPEHI6jSVsrgmX7ZgYkxoH7FGRqn9nBKjnRNon
VDC8EvnBCzLxodc41gltzBRAG7CdataNtAGD3zhEwkF+NR39g5xFc5+y5Wn79z1h
aLg5tfe8pGzE8mE9e9symGYp4z5ventCFiPAU3BWxUdww2ZNyGsIQ/jSA6X6HP4B
4ZEnZOqDS5aQ+wwtEdeJ0CDFea+KQrTJDKN3SawXk2c67r87Igz9RriJsTuLsrLK
X02wPgWuJaKjwuJRnX+phBlnSCzLhP6MeAIT6kdP7Rf7s2Bz7QzM1UEsSsr2p76J
NLT4CsLTK38wR03ORgma0S082tz0wt5w9+wA42dpFPHLKWPW9jjPd6gnT1AU7KW7
lQ85pRZokQ7LSK4JdM/Si3pvFl01DD3tcJSAuYjLHLnEA9ZZmRIeVd3uiBqImt61
9GyMy8tgb6rWEuiYN/KeftOY2ZEkQpA7G8z8Ts5T+oJkFcqvnxNoDJ+kwhL42Wnk
znRP6QlHGo0CeSIKsUjawvjbACf7ouPgXTMj5khefhTLGpCIiUKLEfZlHKdbb9eU
3sum08QTIdZ1ws9pfWBdwdEyjwnqaw0lP24QLOAmifqCK/pJ7bPhKQLBMUbgBv8Z
8FV4dJN4cvv8tGfQdf4xgGraUhScnExEqZC/Hvae/Ihw2YNDDqxC/pib8VfJewD3
yNXsQBYwEU9PauvCARssZ6vMTa98Hs7qJm6FZesTT2QAwsgSC+gJTCQZ601qya9V
gg9//iVnOk5NuZRWOD9uHXB9v1QLSHQ5K5kBgQhJbWeYTNgVi7MFsp1wQqPhDnsI
yNhBCupmkRP4sapSdEEvL5+v7ajyouRrAbN6Dh2BPZt/pyiIYbAuK0Znza08x5IS
HZTtM6izbaSp/F2WVT6EYUOTpmmnNxG/4jkZ34mXCuB+RBzRWeS8J6AbTlSOyBZR
7D3uuaE3jiZVXIpDJ2uypS7qXCHx8mOvUHRTkaCaOAYqufa4Mf5g8AxQCPSf8NYt
RTWtuX3Wkdzk90HFOFtIStljtzgU0RdHxeJFalRZN3AYbm9HCbxKXGZJ7mLbRj3M
UBB1gfeKY53cIkRoflRapnjeBEdvsugoOK65z4U/yxgfLM4XW/LO/xDWKEKAQYoy
84JxfQdGiBiw4BGJVD9EaGl9Cdz1D6h8XqoPmz5ERoMrnrjyWjDU9/f8RomOpqkp
zhXClQBXf43/sR9gtwfYrsTxGL8jSdwBQZ/im7GS+2ZttcPkRtmEI2plgqPIDUIq
azY1LVO+26k48poHqLv32D5y/G2iptHRdtAa0WtU4zsXNItQxxnlrR88CwEP2gK+
iO9sZQ13ITS6OilRBySY6P0/qaFra0T4nimdaey4fzZKk1ABvdOvrntqBTlbwvLA
e6eOvX98u3ImFMgKJRKn72Ocaf3MB3rGi9XWczyjch7eZ8M6dY2Ekmu4nde5QgFD
G2HZLFEBL24ycRL/kIRaSj4r+HVEnnTYAl6/3PrD/m4D/tg64v72GB7AYUMrqALO
txncHla9jPWciEgvPCQuxG3n+jH1LicnmIYC0hoTFTJxwwBMBiwBzBJKIBhjMY7A
oqf5OCycJROanG//MXwVh1WfleF+bAbng+nKcKFoIAF3R5JfOBxuyuB519o2bDvX
RQmcPOL6NAkAgFojcMd0gTT4ZjDfoe3g9DyUD3iJFcN9RVO8ai9v0VLbWbEc7+a1
LWqLAj8ctUx3Q0Vs3d/8MtyqQZDM8npNS7vATL0WdW/XpcPjuR6vq0CVQPyFS5Sq
bNQQ6sb/6tMLLlntwNcQSkEmzRGKg0cIaweatT1vGtZtiUG3RjoPBsiSJjbrlTIA
OAVdyria47IiTSTg/gH8nQQlhO/zf/wotv2+AyDG2LzZYpXsYYm4IL3dwgW6N/IV
rRN+irjPJwuiKQTT6/a+hwlWxMD5YeNFT3jcIYIi0BL7dbgAhDK5iZh+O6vfZS0S
7B+dFGoiScZ/DFmzJxwm3wzaptBlcKS19PjTy4QsZeHYAedPKZgzlhf6gVrTumBu
p6es6hDn9OQ6M1xhZAJnnXAugv4SoEkQ/GFz9Le3RTe7aqTiW+v1SMdmzUOKI9R2
Yxf84IF8p1tRv7BcYKlUiM3VUMxv4DwmkwroNreAj8OHa3noHEf03LCOxQ3I0KdO
9dnmcAWXUfVTc7MHhCpwcgLNQj5SxOYhMakAtyNWSnIB4UMCJ5jnQxEUMdWNct3p
h+ySxMYq3jNxoygUhPbp+kIxa/fD72vALaTQXv1ui8LDpfrN+JGweiT2WmxKGjEy
R6+7M04Lrpp3kSAXxEZuDZdcd83nPaTKANee5oD6n5T7O3MkZFAxN12/7J3wbj0f
7ckn65dZbAELt0laz6jkDRPLpyQ5s/bmqa1Wvneymp+vyho0PLXBxdkdCsFZK2lt
PlbViWvXcO+3ZPwJExsyuJSfFYBABFJPt+AGGSBsqrkngl5dlyYVkP5GEaiTikwN
1msI3FhY+m81pkTHGSPFTsBjXnQ7s5YszhgG/I+tKkaRlnX6oAp9ZabNvkDvN8wk
4D/Nsy1yU/7hpuv8UlJKwqep0QgC3o3Lzh+YuDT0ZhPF7/ZsnXtEWYCx2tDtlL58
xH8MB8ktePsU8f+BiM9kRCLwiVQ3I0IR+Ri/okSYSYkmUQ0Ib9lFIMVFqq2K/Y79
aRIjZp23/gEU+lLY08zjs1C1r1xxyhCHefhPXchM67CsW76uJt9qnvYbHAt7O8Sw
og2jpKTSVjOTKAk6Z6Ukweg2ZGqM5gbSQkKm+8/TN2Dqywh7D+5mlXz/juYzokYm
FynPlhesbkQabUpIUhcIdzY6HUto1JSpWEVPTBJh+M/SNPZ/r4Ds/GaKS4poYinG
wPAwf6CEryHjoFXnkI/P2xyWh1gLjzNjki7hbbGhcEZd0HAKeNvuJGJ+J8berXEP
cCkUYRvexINCqCXgV/KGhcqRYGwS9tz0uyQHaExBSQzw/EJcWyNDQJI1IZGquzcs
g82CSmKvrWoYHg47+sEPH5mxYK6nUuX7FH2mHX3jmKuhRjoLdEiTq5Xeyo92Gn8k
XYITu7mQ2Q4LTC/Qg3IdCnYac1KoeqafmhNvliu4G2Kou8xW1f1/YDQsvBFIPvkP
NHVA2xKnTekTX6mwifIhLeKOC17AOedlGnyvH4cx3A928wI4MhAWuUGWqU6hWV7x
caqC7a8Ed3BZ+71F6uP4MEzAXL6flrSRs+Roau5i3PwDho2hezDF4sTr7oDXVfwx
zHgjHLPez8CKYX9xxtH32uh0vNGjEm15ORWlfZXQ+wROVpEB/cASNkFDFEViBBC/
+MgMyVSFqj3oDtU/Osdym860Ur2yWRUraaINbVfp1LTAd0VI6l5f7daeU33OIx3R
jcZKWWA1isnT7zWZ0Qkuzme1UbtS6aKKoRRyoB2o65/hQ0S7sAGhjVFPBocUfEKe
LnbJhelJtMyqbBgCG5iMBq2ZiwVrRB4JoYXvXAuvaM8bC8Dw/CbKl4CsCd4RlRG9
+D2Is0kvrBnb4mSosVWTCUL7PrrHBbfwpwYcn1pDJOWMNDmJrAX8SrjCCO/dEiOM
eDWp30uoPK8wO3RGh0fmOeHcdAVDu0mNU0m/6BReC92KpFC1h06NVMI/t5oKqwah
xgwMLFmB6u0VoFdIzgrFMCjWRGukQoSVsoKQg5poNiJtyET2C/tOB2/yG/bWvMbs
M3yQBjBmfi97VIETJdHPsr3YXiVxK2x4Yn25qcmSyw3eHah1g01uHyPEVGgvncjW
RxU8SyQ8qzm/ar/qFqal8U2J2KHGE9weYt9SSNKWHJL2/8b9g1fyQjqabEFIqmLf
iAR1HRGkHU8G77aAz5G+5SJUUupy1dyCq6/cF3HMKao+XhNFof0Dkn7Ld4GLPpoe
HzBxfiOx7GDH0/vzVc5alWLFWUqykkuxgrdWE/btv5Me+NZEzKpO34AFwleC1VKr
FkshcQdQCVbo/j3F21kHvBi9N4E3Ggl4AUg6HQp7WsOK4L2t+ax/RdkbjcKxBum3
dP4KL0VoI7z6P6Co+ljxfDPvWcKYNL2H8CNh5ePKDqC58UC5fh0b9C4ujzD/cl4p
Djb/bXaOQZmEaykVwEbqT7Xw6yGE+0ay7xBf4z3h3NOzw50Wk5Fca0uFlRmp7T32
P8U+M4QPJXPwEpI9osH4ZAmDcQQInUcgpzfwk9DW6QKaZuxcB5mXN4z6tjveCS8j
suYxdkl7lcWXpHwtM+8tkq04M6kVtCiDWRKxcyDoOFazqmB4WWxFqHo3qnrsG0Do
DcVFC2WLxsqCVrD+V5+GjmSDGsk9OQFlXUezMR0YhOWh6lHMOIAr7Nq+L985k2Ez
kXKJnyuQQpnTrjH3zZPUiE7XWTWJaQ14huxRDvG/ahfJsHAQj6IB4qY8kjKkY55x
zi74EpEvJzuacfADxBoKyevCYMiTTdOfWO223jKD4CE9kl+aC2SsIQBG06uD4h5M
OTe2U3sMT0xxsuolo78xmwJZ7UUR7nOZugUH8JZ+WHjao2oC5A6JAYJLyjjGUDQi
pKPWRx6FpsVLsWU60dA43mLa2KF3W7zQk7+IuTvCdyj7ho5gyt7/Sqr+c3ZCw1mb
zo0I1tjGQ1UYou8p/Z88lKa6M306lnaRwhmXo+ZjoWFSaJV3CTUWQ2LR8VpMoL1d
kXf/TWEEZM7L1PwmEzTrmnE99J05urf15+xThzLDBrgJ6BSPL/O9mVe2iL02c5c1
LmtyI5gEjlKX9dBzDMAnUfPGn6z9LkgxIQWfVdbn3TSEr4v7K3f+B4dAJ/4eAjui
m2RzcyEpwfm8pX4LVCcvwitwLpH0a47Gx5xlke/XmAhm+2aJ8u/kz5az50YNWj3a
XojT4Qg2k12EJXCMpwxbZBJARfu2d1GWG1yze1nuOhfGDu0omubRpcrPGRxi4il6
iI0dKhdNJBApAeQTUBdfn36eJUV2T++C1b82cLUe5cWi9iZZX5aaPefG4OLHEjbP
SDJiedXIbMgmaMZBC0wOuyUyjy8MDKpsQ7DKPFyP7qMptRLvWmVjnjkUWkleL52G
IawliYF0HR9XszLyY44ETHHonKMMtpZryZ4NQQLX/CJsCWvBbQBcCcmNM/xL2pIO
9WAbseaxiDXCwpnQf3tT07xzLE4VLMA76OeDA1K5eBx3/82nq6uNcDTQHHqH93rj
lmX4/xJw6A9vEshxBB/YTbIe60H1V/DWV2c/+W7ttS3ovUoxkrHGoB6vB0D7D9S4
LNF/catX29zD7/zX4aNUkjkVd+G2zcKpjBTyyh4UMu6+E0T6xrfo3hq4iEQsKj6h
eQ7RYDHdedUw3VALQGK8WxqMp2yFbYkq4Ra0pdbwwKGSvgbwTHACusKCBIrRuXay
cZS6WKcffJTQg7hafFK1KrB2xrixqK6i+6Rx6duSKqUUk1l/67cWMdNodRF2bR3X
3458wBKtaICvAihnlAcRI4536pcHeUEatYo3fq1T6JDellH/xb7JzeWxrkjl89w7
hBIrLYVK4I1l/7AjkkTL4v1B8kGvdBbnhTxgBVlR3z/6KDU6QF6KaArXGYsr02zT
Bz86DTv46dkUTPpvgzWuf7NVl8Kk2xXyQOgWWKrCcExqguI1aGCK93heIYEvNzm2
yN2auOAXBtpboLYJuS5MhHQ2tEUK3wBY0DqqEuBrCTLPgwpKCiOvcpOfStUfdri2
QDwN5IhiwXtG85HHIQAWeeMbKycqVhW2KvmzZjcFZ2x3v7Kfff7lWBEKEkGpTo+9
V1IvhsQxEbh7FRVd1BUcNw/YFFfuFhvn/1VrZ8iCboV38wiTvOPRRYM/rU/dn+QY
Wzf1hc3pVmnZgAEWTrlUurbbtPd32EhVhbiruVn0XCcpKiA03mpWkIgEvyxi8Z/H
bGIMfdLMF6Di9mDlNzvljiRQikhKGuhE8qy5f0w/t9ty6eoZzPS8vNE+k0yhDsma
pG+M0Wytu16esVXUy7jA73Nfga4Bcg/D461Ui10B0/Km6YDO9eQbP5fZPrs6ijHC
YFbSDKqMG6SDGGRprGK7L4XG6D8QFIKCdKxIwDCIP60vE3k+Eq1FpAMKKm8cAqSF
zTj0Auj+PJkqobivGxuZuKjQMaS0FmrzhQUxrxs1/1Z/BWZPq45FOn8lAksAuO4s
XgksYn+D3nZ/4fyjf3673FKV8x4hy3JjNk16xS8kv+lomVGUJh4YPzVyTLvYsl8r
rUfxRu9vkXaXcxGED2IOq5P4GCxEJ1+bStkaDslEHMu2EW4+jE4/cCieTvj14Bbm
Rk7iw15ii1nwt+T4QdkXZpcud16KUtiw87qr+uTZDBDaG2dtu1esyRAxPsOOBFwG
owErGXzq+EIprk0vwXE8+J8JrxCzq7qD7aPihxI6wzhRPT49B/HQkeQqJq0jrjq5
ZX2XhjGSttpde4ozaz3cmFMDD8C1UBMIXCCoi14Y5QsPrt+XmTRQy48Ft5xrnyHK
W0INvGBlc4QMKjpp/r8rxpKAP7Q45lQM/YI78Woss8I+RUTxvtdYi4/Wz2LK2Yn/
KW2M8Ejr/AhB+JZVwtaf8DLhlGXLkWodh/ghkh/kTMbgOMWnHMW1CEbn4z9Q/pKH
gldJK8JwqBbnnhx68Mah3M/v1H4brKeKPMQ8mUCdE6JJpBPgc8+kuKQ7ls7qWLEm
jS9wX+6SHZVHymyaGm2ws4VJwpuZtMg7jxWunksP61dd8AU0gaNeDbsCku4eZ9cW
n+4P6spzYznDtpxcLsCru4IiTX5lXwJex5AuhSFDVQjYyUG+Lemp+qYyUdmnqp4P
G5jjCSWeGnHdBj5yTB3F5GK4qBZVUT96NFIH0UXLPkLhUgl4QNGNLu2a6n3Tqhcz
LnKOjhZJNZZ1eH3LSSoWjaD2WW/jUPIk5Jl9nsMT951I9807Ai264eCwF/iujV2O
RZ3IwTD5MUDQZOXFqLPBgrmRna48b4Phl56zVzQ+kuEVv+7DvkZYUl4HqdUCYnEp
sWnvrP0ZnJVbVZX8Qj4GydxPTU2CQ41G7LEbWWUO39AUJMcz1Y/xgRGsRrsu5MXO
8oxBHcsi9AD2Jt1SPmwHnQo4+hysybep7Ks0sPp7Vjjed1vYHZ1nzEe3kBVjmUWS
Fue55u4kb/HCoRneb8va/pROjChlO2c+1LT+s1A8oC/Q7xoiql3eA5aAJd8+eXMT
gsZXZu/ncHPI4VUhkgAITCBb7HFrmKNbk8aRjMB8Zm8tCjdhs9MEaKhCdwTm8tA9
31ZMw7/GCCxu3+b6bg0hsyoHg2ihcxrRM13EttkvNZ1DqtFy2MHRtFvIb9LoGRG1
mDstfWVxxOMjra480EIrSd93sTRmCsiRWgFp5ephRKIpH3RObIyiMZyV4wSTWFeM
x0Z9ScyD0sDCqN5TQk+aj7+6+FoHjjaXu09Iq86tlfo53joLBiU2huI0/1qUMixd
3tlO1pd5EzRwAmyDgnPM+hQ1knB2iLzf+CGOgN3JR77XDEsp9hF1geQz3EhhcNBu
yW1V0I/lfumPvHNxooRujGoUaecKARAFXc1xvfX39asxH1cfuNT9jj6H48QWgPhL
KtKnGGSHzSym503rgZfL5W11GYD7LfTcWRRALnZGS/R1bMNZ173C9seN2b+54CMF
h+refWyKz3S+ktk8N+aTjGZ77mzlVQrl4bblE1KVVhoeCc5a5qcwYvqjl9VVqw6t
uxKOtyTdhWiEXW1DBxE92TrTSGurUOkJk3oc+Hi77DuOFQRTcva2pf4FQcB/yXZT
VFa5DnQlLA/3kw99e/7YtlKGeQ4767XLiofhWf+r5e8Wfwe7ENF4C7GwMN4DK56B
I26ss+fRBTbZ2OtpU6r/xhz+VKsip04WvmHyulIQH8+wQskieGuX+cQPz4emn9bI
kuuwUfz50v3we3AZSkrWrsM0SpTh4V/oUBHl2Oj/6/68DO9ErwC13cmh/4+I82Vu
kHOA11Nf+zHDAPE8tcoR5YGvTUz/KLwuZhKLV4NVsU2NlAvgZn1dWB6s9KKVzg4N
8BaGJvSfFkPBdR2Juq5RT9IUxFoHkYo7sWmVCDbIndcEfnNxhFTuTk8SNBQbMGFP
1YSG08DH9eIIgfAqfxovDmesPZzOZyr/CwgKhDuNOtVLyorhqlS049leCVkf8iBM
elc5AaqcMmJBINdMbCdbRZK3rwYVD+y5WzPwoMCfW5bdk5HvAk5JE0Aqh6oPsdyS
4zNksMIqWDm7bUF/6vWkuD1uTUgy9ZCjcHIcKbl4CIrepsMJJslvrP+Z7ChvCh1V
s4PeEpAtqf9UtUU+3xNu9b7VzlPZcv3Qdck06PCaoa8o/xnNPuZhVZJac4Jd6t4g
4OHP6A035DK2x1+OX8IOqp2ohyVZne1J/9B+Aaafi/AWWPUQ+EgnErSQvWzfqgHs
UlfFHRhU3Oz4FFHCPKPKM8K3vWN2Zy0z5T4LaowVgGp4KDu/wVjSKp6CbecygKe2
DpfSw/CX5yejrzQeZG0V2UwsKfTpgNpONagTxgpZLfFxOv39OxmIDQDgcZr+Wutw
WT6k0Er+v9zcnmAsgjmIq17FWeT1qSpYDCD+ZiaGtxCrGiV5+Yospw1BhCBxUQpA
FW3aCo4qmeVMxeuqchHaLVc0H9w9A4BorjKsNFlEMwATpK2pWRrsKTYM/fLyWChF
UdOicCJJu7tP1cyjaIlX3RBAtDMEtPSIW2RgEPuL756rrNaNz2tgaqwnW77k6baf
g04f9E/U1BYVrXCr9jZky5Up3/jpJV+b9dXkDH8czXwCrfdBtpkJJzTcOTjALN6/
HDLA0kubDowgtrPS7H9zc0qjva9UNt1/Jl4sCqGPE5MfXsYlnE64Yjp3bo3pxCTl
5ajNy19rek/v9OmvqIukuGUv9hNCy+WyrvNzd8RMWWW8PMooO5EP65k45Mjxu6Wz
/qH3/Kg9VpCg7l2Oc4R0+pGGJu6WsYbE96xN85SAoglV5rMFG9L1XUY7gsjWKQMp
RLteV6FmEQx398geOvN/iwGpFu9AYLlerbA/PDh2IjsJ26pZsQVlSG4ToVWNfXlx
L23GMya8uGyQ0raJqwUrLBTU/wmtYz24rfYj6OHd/kaqzGzHP3R6PwVUDh8/zpjK
anGHHB8IeOQ/ayOz0BAKXFPYKoUVEEVrSjnV4bYcQbdHKB5jkAP31AEaXwWxlbPg
Eix75EaX8lsVWmY1JeNwNaNNS+1YiBACAIjp/CtIdk7xvoSj9bgzSccFR+qPnXL6
ib9NNQq7JV4RZXMiqO/rUfiyt6a3oOXxDkWrCZRBBz0Ao9FzGnc6ABYndcKLFyO3
m/NwyLrf87eQOX6r9LiIO3hlkiQt/2hB7UE4P8ozqL8QRJr+GwOvDORSUkfkbybn
2GfdZTuly1gBZB0Z4cJZMNeJaL02ItJpwhcFLxMIRO8SDkdfe7P4VviVeyFli8bA
W3yDDoDCcYrcjLpTVwxf5DtGrgV31WQaySHi70RPf0EPHVs7xAItkrS99aWkp37+
uMHdxWmdR7J5vTpJKaxcj7rsnsjqm8xruoRBzU9QN+carU4Lm/LRMYU2ri7j6jex
IMzTSRctPbqq3ZDehNx5qyEJYdFwbkETKG4d56ikUb4BG3z7OL98ngInQkwCIhIw
Ss5dd0Krwf3w7jdDlcxVtLpWeV4LkAGMHNLkbYa01X92CTqlL0BsNc79HtrwcJVy
ldIc/Mhn1CHbFPsd+hsRsJ58aCWStALkxjiYuN+IT84ejBovRf74v92S0ECNjhN7
jHORGLdWeIh6U858i25FqMSQhxxYOBnpvz9z4ljCZCiLA0J7orviXk89MWyN3jr3
1iDJwneKEynfyVqhhSDLUhONjcHV6K77zLufeW1ZuoChG+3BNQibEO1HiHSeweOS
qNxrv/ULezh/+qeuRz+Uggjgys15AwsBXAUuuXFGCZ2Tue9+L87subC3aJ4whX4b
ORM7KneDhGk8Qhq9wMyKzR9gEt61uCoRtE4DNBxHSrrOfEoIeIjLPp95hjqBR+Tv
CyFI2IvidZR/OYjGYipeqzhvEmz1wOr180n1A0/sy7LYq6cjvI+L84oBZIkBEM2x
LoDD752rVsuEaYXDeI7w2zcTIDJtTFqmvK1NGasqfT6Uat9RJtEOsa1iuelN9UoD
qxffDQeo6epvSGCvQFYDg30cXpeRwWnolNnmw/rePXPxZB30rHG2Q4ZdovxR+8Bq
x0w7S4JGYMma4Eqcq+HLxeF6Fj/mNhMtQbp1kLf4S0vvgzprvr+mYFCozMrJDLoa
oI4iZAQKbcoKXlT3E18BVjvO2YOgXHLX8QonYuL4+EP3AmZv9f3o498n5vLCYQMP
aZv3lsnC8iKAM3pzesb44zPI9hVSn0FbSiGl9iCOQZCnj0hlkQgGD7eqbfAmcFHJ
VygkuVGXrsCONr5Tor+UT+qy9LewbB3Scs4X13OeqFGf62c6+qfC87flSE2H80lI
6xn4I7QLAlU0NZogFDf9BVCzC1S40GNCnfWFPQahi5CJ7sgoxtnO9LSEYbs83xPZ
LH90ircMC1w6Q6AY+h1Mv2W0Lniz3WiTiOtaoOTk4G9HRWF6u7qp1F9gRC0kXBTd
45kPXkSW+Z3XltBLb/Gmpb9H0zIjKuc4m1htbWxc4fBTo0AIX4niNI3jEqhqLBiP
1Lzj9BqIyHWTA8Psag1vi4EjXoUbN7T6IGhlJmDFherql4dg0Z3E3K+ngmOzf8gd
kpwrYfjYopm679IFP1atJjMRWS4iCrPV/Sve6wZMRtGZsi/2bN+Rs4urJOTfdR2Q
yG642mdCSWKtvf29Q2qCt3RcFhrmT9HobmrBG/QhjwjSe9bQsOv4hBeDVslH2EZW
CpdV4/LPRYx/HSGFHLBg0Kx2QTXCHP06m0KX1u2dQpbAW6pKWrEq9aFgBsNsYHa0
ytfuBIGFlIdITSEBERQqxPIwG+WkmO1mjn8lwPowalWwrbD+jYUUowlwatj4EeP6
q6P/KTS/5CYqx1NimCdueT/YkysgK3kugvBilo2RwiON2ARoLvgqcK64w+nOXIto
tZeMZICOgYK3OTVz4dVy8ofBIXI2tWxktUpZWbvF+SpDPgYjus9hrLZ8b7z6Fr6U
YwsoRvbG40bJLuM3cW7ihpj/e54hN9/sOT2JfXQvLpnRD1WNVrnSXbXFDdJyxoe3
VIE0vlMjtSwDbQ2EWUpPU+lTd++gF7XVEhmY4NbNzexfGkJNp7fsRoXjO8FBv0PL
7/138sROrWJB6SCCI3uESNBz5dZJlQB634domd//Mp+KQWRy+UR7qaUH2krFnQvD
YpHSpfy3Hi97/8coI1zE71uoj/rWuCooyewYELciPjgTxcF0b39WIPtptx2kgr4v
TIZDHAeNQNB22Fji/1DjzdEo/uv/069jlc5Mb4UG9ND+YBgM6z6mmpLUoqhYaSqV
9Ynjsru52FACCLm7BsNVCBftBMfBpEMQPcT38hjGt6LKyCuPhmlIU5QEXENAtYzl
glNs/V2myKWiRUkd9qlTatq3kn3KwBkYSa6GMwvKLiG5CT3++yg6WfFWcvbrC6Hc
oC9KpUr9iWStUi9MvjGbbf8ic9dAATHUKYy4gEnDDzTRBxI/MCZN25OFq9E5eYqj
MWGU27xUhx2/lIvpxopBLvP0A6lF4gVDswHS5bPhDdYLDv+ThVWNDWfI6l9tXVOw
f+nWCRpDXWTJbOijS8nR9DN4gAnbpl9g7WYwLeKot0zTDxJDplG92Ynltu+m7sGn
s5/weRBVw1M+CJ8uDBIwEZzBSVSUtZwiEIU1dCdK+fpbUUgOB78YJaLWJpqlAW7N
I+Nib4c2BHN3yWQuPqi9QC2HR4S/olbeEnmRqiHOf0XMM6CMsilcuT28/Fa/94pM
230KyJrZM9QzC9rpVtUTOJZVN7vTDqknlAQCzrHfkHbZR39yQZMZeK/wiOUGdbyt
KB+26Vbu0sFl5OVsLXBZGf+lEiw+YQ8W2zhEqX7SaOjzoAlOOW8xx1snKZxHe/nQ
/KRScj5i18QvF7ZEdjt75r2ZgmtBH8wFq0yLWNJiVPCX0joYCPPBKWiGeybp4VEd
8fTIhz74PMuL9OKFa88zeEnA3VSznOgy/fcvVZ2o2yxENM/I4GUx6e8kRW/WeoLT
IydRfOKvMqAnAjUmeZx1Bm3hlNZq6AxYt7QIOO9l2kvsMtW3M6JHHLcZ2C5fSo/v
speCQm5KbNwUgmczlHRs3fjswwyheoozuMLXcs7UimnLkhKYSsicp/8mgw5J2gnv
/eH9D2T9godP7Ap9tIlEcbcf/c/8AV7Iul6QNiYeeEK/ICJJBoj49bhlTjuAOq6G
B441sGeskdbQh57gQyiqs+nJr315IQQwrGEYQOlN9kS/hSV2PwM4p5UaYgilqWlo
lR358ECr6MR+f54JIIUwD3NnyjqQduirO9h8i11rd4paWrUFM7a5FiQ1nWJ7IsEU
mPaM1IoTPs+WAqe0WKxmMVi+POV+KD86ELa9Y9ZbtORN42jVhZ+19kqER3+6t0/8
p1h3E08f/27MXW+L/pQD4Odlr5QU4T7kJx1LGDGrmDk8s2OtqjGY0PzMhXXdsIQs
hzt0kKDFoFh8Po3R8FuauJ8zvJljhWKeyIWFGDNw6UvW9UgSZSu6heZilTbmgrUl
SOF8rKsqUo582XLS/S9J/oYWY7WaBMtz5QIQZGsqWXeIYgffSrc1LZ7ThMM80KPD
XqYS/vTbKsz6A/9IDi1/wfD60KgJcofZ9aNaR9QCaF8tMgexJEtStWQn52nJx9VL
L0eYOYsYRFPLykoZuxOauQp+O6PI583WQSatCvQo8RfPgtB7noiPvV3bqEmWX4bL
uSyev0UvBuxCb9koBy/tuRhvQw9srkJ67bre+BATYpCLOYQ8y1cGm1iyzDz8zgv2
4pie9+XhVF2irpF+nblBs1g8F1CBq8reQuydNV18kK2AJ9n93o04MwAGQ0Ic6G9r
DnGx/eySdQjBB+UrBwMywGO7WYFR2lcCtTUc0wZF8oWtZdRHEFrW/7CHodKrjYCa
1DkJvGpAMQcXx2F93AX7mVYWJ935WOMIRWis0BFY6Y6iNuCnE4juxMgdZtH1nzYF
2N0ea++FvR14PmsWEWHvUyE75FRrI4LJyIRNz0fIyzIO0SakPqYnGO+F+BB3JZ3V
urpWaKEfXVQp6eHb4jHhoGpWRl51xb780oVJ3nx8u6yHy7jnSNUH0JP03Rp/v+Ev
QrwUW326rVCJVEShppNhy8gmIsrn2U7J5O7ummha0sGm4wVvrw/6FOPUZZ8Yy0N/
5Mu9fQcu8IF4wzFmQnAiy6kb0ZQFDD6F9f6k6o+72dwE2ByDCcKkYsX3WuqLd72B
KyWUmdcC6AReOR5n8z57Vyv3x1iKs1o5V3dFKyINDHWL8MNjL/DduuNKasXPUbEb
LIwR4Y4p2Z3fuvnt2nT9RvDoUEvd+v7TKLn9YB5FFZjkBDJwUx85F6gPd6+u/eCq
vlAaiV0/lf2D20t81fAJDN6pFsvpTFKkYMIYb3qBvVkUw7aPu+5d4HjVTy+vZ+oN
6uZVKZmab+M+Grk55Ln7ggoC3lfQHgYJS4dhUM2q+syRzKybXMz6qXgh2ksH9gab
TvyAeP4rwfbxug6PnjoUNXtEiZVzwHSQJ8kUS8zy7TFJ0og/WwNQlli2i50cP2O/
th3iGNo/r2e+gZLBNYQLQ4NQI1geFEz/8xqt99b86ckn5YRo8zVn6eI72w9Daqjc
TeORgE5y8nPwfMRqLu1zaLFdelcdv0hrKB4Zq/HmiLE4/YeaUqIZYi1rkm/NRpkS
htBwcE1dTeZ7But+Cv7+u8zXnWdiu9XIczSlaiySIPDyHfid+26+FKugbjYKKGdg
wE7EkS3q12ZG/+RgxokFox5w2peiZDaiZ6h48DzLGZtdxvnoCsoLtVHk6pSv+93W
IMSG840oro6PK0fOLNxetQg9hdhA11mQwQqw+d9fTmNZ5nitktYrfvBu9Cbf29nK
BINNOuAlWexYtOZmAQtN8ZK3cEXbrQkd+FpREGaOJ0RMiFmXa+WsgyCosSH0jfX9
r8JdPREbe3cYcxkdqjeITPqJuxlKTPVrh3pfE1m/zaRnm80vf68Du8xvgTghPws2
BAarr9paRgLuNpAvzvVT80MSugpGJOzbVc3e3Kp7ukPpg/6q9SCLhk9BVgRs4Zw7
KztONfyYWq50NNd0qzpu/0VemP1A9RXKyyLSCC0/Obrte8SpXo04xC/lGKh740Ua
fYbCEMJwbM4IX6QzTYpQbYIuJIFCsIK9YMSmvw73mf9+gVmXt3E1qmC+o09IMmQi
/0uOceb4uyM1IcR/ZEix4/ngqgsDFrkb5f4MOj/uFWh0Z4f1ACemg6XB7lzixPa9
iKMFARuu+3OiVapuSxEn8CIBdJM6ISqdMhNudN+0fQZ5nINC/sMg8NPnFxLkXrj4
ywADQENbKWKXNCgG7H1x2kG6Iy+h5g27vkPwcjrFZVAHF0zpkCVeaHTdhJ+H4+cY
OO9zq9LVtwSTS3TKoFu3MZZhNJvbVLC8xsjcBoxNQq5SfuLstYYFaLCEvvxxMGjZ
oIw5HN/Rvy3I3aTr39HWNTO2W4Gc2dXmg+m6f3tHpzdl1nsh7Z/c6hzXH6KDHcsD
p9AWjf/Rrq88GSimRfkc0xtnd1FV1OrKu/6xN4Uki3DIJYaYMsxkRmO7cEuf/w/w
AjZjD+/dHtfbTvgnGRey7CCuapS71oZZ11G8OF7rcHAYUAdaDLT8HdlCdTcWEYQi
7Rhc6ouLXOxDYg5+BxZKsKJ3vJrErv62r5Tt+baGLgK6i//T/Ojqr668P1oHCfLP
S9sBbYC8eSd3maZfbL8E90Cv7r8x8AaF0zwbkE26u+7893OBPqy+uXsPUb0RsSNW
cckCyvLd4kDdIvXdcxKgOXMg9j6Fruy097tbWO4MrhPZTiicvt2E15HpZJ2pB+eK
FmgT42ejTBkkitWvklNnmv1/qpNCECqHIJLnVGiGj12OU0qgtLvLv3W1egR97ho+
6CDHKf11r1yc3arjFaJC/FJrm1FmmY+FJgtdfnP5fnIJShE6iMUpzZh41K1xI1hX
0nv9QexKDULLNQVmbFBXC5RevldcpxiUu/vHfJLwBM3tv1lmpsme6PpBbxtkhklX
IweWMQlk9B69XQnU7VCjq3Pj5OHn9dC45Cz5cyz2QRkYcx+pu4S8AWidhXdjpBez
9Q2/78X+li5Hr8wKbErrAeRIgNxdvW+cXeJv0ziyX9eU50iITybTA5jmnHKsdxdh
C/AJh9BFpcJungX1zDJXeGSj60+CWt5X8B6F7yKa6PtV946JUX2mxtD5IdhW95vd
q+oGrXafDUPPTTDHr2VDo+ASUTciEEBbC2rIEfjgd1q67TxLxdbeMeI8aOw4wp1+
VN1t3KaCQedpeIlFmG+NAb+1o3m20qTmHlE8AEBqLcH2zyqK2cxL6i7dR2y8XZvF
MCchIgAzMWsgrWM5CDfild/CS6L9A8SASLqNnWw+K7WgLcI08UFzybDGxDbCUf2o
KKElWsALtZyAm0+SRjC8pUfwDrOu+vyGigKHBCk02lI3L+KJfdF64fEWO4SGHlQe
0lokF6sTU4rb/TiQ5X2eqX/FAafDsV3M42CeXPUQ2U+53hsoD+YXBj5Jy2n6HgG/
GOSdacSuyf4SepBwGgqcfn6O/YiA9pie704tPlg0zq8AAgoj6V3q9HU5E+xtpz7e
AXcFR8nw4QC4wmK8qHtJ7IfWMvFCvKgQeKEV49ldB00amihXB2++ynj13oUzlHi1
ARIytGl+4do5MKmR6gWDkvpdk3iqtC+GHa8o2fG86BUEq6upgbznAMV1YrYLXC/H
JgJWX/hS+YTi+nmsCXwuxUJkUyg51rO9LZuw2Qv+1EpRknD5wlK3EF72DMD4vUXi
MF/1O6/igWzKChw0rPR5S+uTYVhqrz2JrdyappH1uWVw3oHRukNWiFkHCWbsgF1Q
U/7/wN1z5b8JyIyWLoI+HLmpl4lpckFeRwMRwf9iZ9JLSe2KLpSWOIePko/f579S
e6T5eyiLxgOiH9BeLIhUzZA2pkTR06r4UR3jRbBMBQobcS8KKrhHNpoXClXzAOqm
VwAQzZtknhDTdZfHpHTzO7MhDYhPsFQfU2xRtV0F5e88klWTDknINQKMsb99Lr1B
rM3S9tRHhZKQQQji4uak18yUOFkUoV3ejPUocLxWOueID/lzayv7/Vrrc+wafNww
6uuA/9WIE0HiMyFVH6fTsyh1MtIeS99uAdovslV6TCW4qPqYjmzxh5oQUCQ+9o5Z
JpboABjLTOps/O8rb6UL3GXBxtqksTMUO2XLRoURFOtVPT18PX2nvN0n6KOQ7/OD
Q3grCmjz9DRzM18hdnfNaeGQ4Z4MwvS5XgUJJ78O/+NUL6xyHezPTgqMtw27yoWW
VzPgOt128s82jx6aaDkj0yczjqBOERsC28OUb8AkNLAZITOmcJ62jEGwb8XTADH/
+VAK2aKAEjnC0TafTq1gs+INz502df4x15Ti8ZlUoKrprRgk9aZCDDq4YgHH2b5N
flW2dZodPCRv0abyUczniLtLqBQhYqT0PjZv9AGQ4PpaPINhf+VLhHNgCXWSNOo3
fUIf9bH++POYG+6JC+tit/sMro+FAhilu1Gf3JdS5asMXlhVOEjSgLQ50MKGx9ps
vXj50dSjVef0j3FkeOk+Tfki5OdsHtifLS5+NT+kgrkeG7mXMlxzmu7VZBGWvVQf
Jsx5uvvHuL4qSkUwLPmnklpVy00z/YUbsh/4uGw/KOyE4DKmUOhMHdJD1r/uqpe0
6c5T/r1noQk1x+WxyfM/K+A+08gPsCepyj4blpa8XxkAFn6Dj+X8QBxn9DXaC+XC
CSQShNGGteCf7s6Nt1nh0EI1NbkVXfULRTSYje71RFlxLQlkVEWUvqsWX34iqPqc
EZdYKFJ7jhMjtqyC8lVUsIuNKBm/s6oayECW3pkbHVlRX0XebBqYnSKjMdC4bATf
4GF8Yff6RI/wbyzqZIWx9qiM8LMgp8DxZf/sWENbTQd3K/zUqpGBiAsjQgbcHlg4
rskOGqUxrB8HswXOA2yVbx41brwI98I7s8JoRh3o7XFTTcd7oH8rwFSvQpk1Xk4D
fvKVXL+YSzIZ0pT4R6IKLtxCeFpgorrtfDBfyKfBWuiTy3a7OebnijkW3G/O/nsa
iwwBx8meiurOYu/GxmueeYs9dIZkFhIX87qotCBLODs8hlkxfSzWcYewfkMhQzsF
0p4N4XnVUaNsERTq+lqC/Ie2IsDHuFZLRKmmedBl/Grm67ChIsrbU4nWhBRsrmJ5
Ux+mLysGNeqCkiptp8TxEYg/eAXaEsBzN5YDRROjtvV2A94cuHbWP2ScHFnnJ1Xi
zlsoXRmTwLMTVQNhmfn0KKQWkEM3xyIOU9pevEDqaGgwVRoeXEHEcm7LI2z9NCUF
qEGjfnksHliTujtm1ARQ0pwdIBAtRRbmMZM5rmbn7AprolYQJbLoz6SmuLhfe4rn
vzHqeTLwv/THMD1ULWJfiZiTfKlE54z1oB0GOuad23IZji89toH9hmFNvWuDywzi
3sYpKp6LwrGIu5jWu3mGcFgJ5IQmNrDNplhK1xPWtVUZ2GoAMnZU1cizpgWk3K0q
6k5KRFPLzBPOExdTy/megh3XEYxcpPlkgud2RA5zGyi7GT2kCFflyckLY+XAMZX5
Ggaw62CEqCQp3aTRLxUxIX0QVFxRVnFMoX22IGSR5h1nmGihDi//AKxDyEP+N1Bu
CvAaY2v+fu2yq3ZRr9NXp9YFO40NNwJrkoHUdV0icPR3RhChHnNxspKMvEwVO78g
c/5mH9qby31v4/ITKGogND2Vqa564LjPQ80Y5o/XPBP0vNLn+IdtWEqolEcN4imE
zVwgKZCt37rzsuD09lcD3vCx3DO6N+dfOGckmsb3XzbFKeHbAlv9GTico1v7yaMS
biP7cd+xEzIpY7o/aFToVo9REgJa9arQfKLodwNVkXfsDuZWXXUvVAU9xdLJIKWC
Weg3RPt6PmE9sJOmmhR1ovw8qPvJSZjoq9b59pGt5KtbbFEcKQ3047psjAvN5CYq
dDIkx+5uNf/O1C6509opWbGjhwAGmiBUgcaL+bIQm2ZjVSli/djlZd1Ut2fZORwb
LUV5/6/bnkJwUYO+5MSDvPOZ4nDJV5Lv5JsTb7zJ9VeF9lKO7ldxV9hn4j3PX2XA
qflsLDSXzRBp8THSlyYVWZUHVYTqBMpeOzLgYmJM5AmxJuPpJDDFZS4baBv6BlkY
HSU2TTK0m1ejc1pmEh9S7ZHBnc8rOmlRpQrLxzAZV9RzhNrJJFITWOuR9LgGDh6k
BLoJY9+ACZX8HQ2pNmCaMAL6TuNjg1Jc3zwgu2zgfSu5OoO08SGiuDFXLernIJnD
oNM6bklxMguL1awDnimW/9UfCAKGQY62jITjRc/PCdBkNVeeVdw8vPxCJhOkiqjV
m1+2YvutDLXCJrrycUQ5XJciaeit3ZUCxfhIiLC/wAgHjyelO8pyFhrC5icNFnUD
iqXxP7pnSjqd8vbpY68VOfCyPQTZV3e9Y2aq5PkA0HNu/L9ifmK6wW1Fp4SRsAro
++eFQtnnieX2P33qVkxUKgGvXhn/+/kLYkYhg8+/1EkOKcsw5KqxuSvVpUZv1CN4
yMT+t3rPxlmfNFOHd1QBZaWIC+zPcAryNhzENRSZFbgMjpGR7oMHbLrKBwI9H0uP
tz8bHhzTC/1e6j1Jw1IcXVBRoQlye7fAXbZ0/WXyxjOdzyTz+UkZ4f3XxIWp0MIK
DnFQDUpWPtQ8K4Y3Ma/+kogsI0rKjRYBR5OobmaDMXS4nVsjgoj+76gPzVgozM1J
sMO9C9pNigJizeFVpcZn7jHoE8yw1rA4LPI7jWcdM7KFNt6scwXaUtb32P71NnzU
iPzFdC0tP7Pei+HewZ4CdZErUTyYsdzm5BQLspo/yBbpLMWlb6499U7YICqd7dQA
j2tPRBOC8Eom2XSch+ExQBJ0P8T4FewGZewiSvdaLZJ7IEjanCfQAsrZcEXjMDnN
gcZ5BK8O5LzGx86kOdpB/skpw84QfVLRgpMVYomns5PwmniIlU4tx7LMbhw8GIf8
0bsuMqO3Yth2X/QKtwi+PUnwlZC/WeoIRW92CCaIQ7b6k9XI/fU/TlHF3hTtFOiQ
k1AilHWsG++pf9xxhkpDwhR+32lG8QVXN0lhtWlUCPvRuNDYDDtT51ra0GVEplWo
+cqkps/5YWf1RqxvLbt2hhAKUmvfWxOK/21CsDTckuhpDPDyVGfjTsrcsUbZbJgZ
spT+aF4097AjaCuv1OvT82BGYfm6NJuFB6FYTldyu/LPlLchsBNw5fa9GqdLIG9R
s8/8e4as1znsyAa3JKawhZQgC18Qn1VjoK5n7RDpv6AUp40YZ+C3wvjf86hN3KY+
ZAfIUS4xrSzhjYuOECpsDTyuP6xEi08oNE3dpN76HnOVKCB2GNdE6AhnFM1DVNpw
3BdZxETJ8bi/CtBoSGcT58VOO4h/hXLWnXdkMzJq+1YVOQQ+R/PM/wxotp52ntRT
zONBcyQU/ODQE+PX81HU+3Gmc+HxA1Wfl/3rnClkzoGn0Xq+bGZ122jhOs5vAAwU
CBxylLKNnLIS6mk3ZtVbg+RqVBWYj6vT/OL7wSKW3P0oR2tKMGpm0DLt5mtLqf8Y
3LWt+bbUv197M2Dxh+KTxRqVFA//rn7+Ms75aS4kiaCxYAVBhh63PIJmf/B5JAO+
9auzizWFZ6ekyY8rFdfp9nrLI3d7SxKfG4vlowMsZN8kU9+Fr64msnkFAiClcv6e
1ZTxeXXWQvBc4vjaIesb1+CgJvK6On/8N14lDbG9BRKmIPSRgLyLLlb/arDt5vM9
rFGbVZ4ETo3wBjyjANUxVsF9TP3EAOL7IfdjnVDctmquGDVUQMr2Dxp2XZAD0Z2V
ZXw+SE6/LrnVvbCAPddH35QPE5JXR0LoXAA6CPPksySRsDMq7KxLIwNQkFnSlV/c
EayECusK8SPEUiCLk+OvpUDcoNbLYjfeZcgPvjvuFDvZV9XYzrIgAQhSf3K3gmN4
7gvV4Hze/xfDxOyzCj0IjRYqIozOlSov2U5tTt80zO42bNbJSDeGvGaiPGD66Pys
jOO/K/8nrZIZQHGQm1ZavOXqA/o2rfo3kj9p2s/ybEMkYs4VdIsXL1SZbNZefweB
yKfQGj3Ey72yhMgV0DDiU/l89FF4wBOAvohxwxDASCsKeFHoiRZrKWkdvzQqUcvC
ek9ZJptQXRR4VXRRqwWfTVNmymlsrNXKSHTdX6arRGkrZYnFO24tEmxhwtb9iYEi
YO+OTT2SDYaXkGIG/qExa8F/HzeiY/4gN87M4GeJj7Z/kyZ+cE5rbm8ebCdEjY6R
7Z/xU4/fxPP3BvbHZU9Vr6xMp1ORNG49bZCNgR/8c2vsVQV8nkjgW5o//fTu7n5o
JnCEjCFzN8NDiUXBnAfboBlcvMSjzB0VHhC5I2EZyYm4W01dPAnuiVlorvjuN2LF
S5aHMf8aniZIbg0KC7wdpIOC0pcp8pi/+Lt5XYxzRM5EClO7W/GzUMgcPMpgGw1S
EnoaVp/81/zJG/TKpC1ZZRqkVBlu19MK63RsnmkeG13LjF+R/DCbaRtFJ38+OEoP
envwmSqWlhIbNWJdLe2lyY2qIhX/QNFl57Ogkh00UWei8BI04jQ6dZPZGxCc0lmK
x1WlOqyRRcALvlndLdXvUk3LV793fEUcNgBRsjvELQlruLJaxcgINWLO+Qir3WOD
4PVVy9hRxntvsgZwnMIqtSYrYMNI7/OtZ8pqCxHVf/gc6U7g1oWAPsKKE5LfYfnQ
C8xjwHdw1owc9lgvm9f+/mAV9SHJGi5AFtYaQS9dDEbYvPZcWK7oD1AZ2biR8eE2
wG6wSkKJbZAz5C9s2qXscAeaO7Rs2vAnP55n1Aoky/ccpiZi0Ley43ruNQWMlacK
srDacIvrgvtqzDoYZyUWmZLsnuKUFtLVMYHyOIv7jGF2RbnE3S3Kt4eA5p3e7wqy
/pBFH6q5U8/qwDYLJdC/c2DQCTem8SEbv7WMstMcmRDjRzKSToRt3bNs1MkAubhG
iTez3wICg0lOWPMQvZqlkNog/OR7syye5qkIk1O0tQFda7Nb1c317YedQZYJm9/f
pfL8dUi5xlFd2PDFmpfX4m4oR4wK1Yp/ZQ5S4IY7itNADpWDJ2ZPmkwd41NLi3l8
5+46EAEoJYDfiq31okPWV63lhP06cjPZ4k7IhxJXRoeThOmkMve96E2D8/UxZlap
lcRQipJP2Jb7AQLfhtT5IzalPMSoZNxMZ6AG4xjVekb9g+tjRBTPJd/y4H570oRh
Sa6jZMUhluoTpDvQ3QXP8O1475QgOewo4NL5+xzJPPIgmvrXULSxusr+SgWo0wz7
tC4KuliJAoF9bgCRLRXtMGTf1f8Op2UQprdrIyKGSP5fQLKKyQKuuTftJJRE6Gdc
gvd1SVSTr7v64UAh6Ncpqjww7NMsxdMNJH0Hn7Ng2ZuT5qujXT+4tybK2TkqJcLo
JEEujf77z14CURgZ0jlmkilEtsKTLgHYGVPfSN4I9vjJOPAUvs8OwcS0mwqxo5Rc
01mnZ+Zp2FUCx+ur80lJYpv268+wA0wKJCqSkYjpHKV8gAz1FsWLcpg842aiVP4o
aiEeAk5wVsat/6YMrDa8N0t/sGhYGWeGqBXsdqYM6Zm1GwyeMQmI//o0T2BHMcf8
nJOjTDTl51n2D3JKzk7cl1O7INJoETyEzG9Mrb+e+KNYuWsDhip4pW04i2ycZlsX
qSqazDjEdpqmgzule5jdlXtCGYl8+s4hfDsasZdj653cnsOw4njVNioD/rxAHyEJ
RL+LqDF7frPt+ezXLlf2XoPx1Yg1afZBAAcsu42ixv+JaHujVN6CkPN3PP/iJIvU
E1HJckxKhxy3rWhMK/wYCNyzTMez8tU01n9ElhhERvyY9pDK2tVIpcDFDv4eJTbW
7dxB0ZgqFkZqpSoorsWRljq9ppVEEq0lm8h/9dTMuMJgBPwpZ/vdZYWrC+f0tBZj
o/r3agccButeK6uGG2LnfpTkubUtA69fGjfXFbjw2aJ5CIr7LRg0mlgZEmOOGDT1
9/fC16hiJItx2h0mf3lLy5ziK1PPG4qJdBvCWjegOpiPTK9TQohBFBLCOqV7GpZy
dok2IpJ7VmTEtILal7i/wWIO5h9rJlk/iSwE+xgFYacJiyjWI20cwQVB30tCoDml
mOxqa+IxGNzOZNinxnueFEvtOlo6p1IvCxiyebVPFZ5JNnFk9vdILRIY7b4sXw6i
8tGkp+2c5T6GdcW3dyBqdnIjsqivKzJ+Q3pvYdJfMhPz2H45YArY5v9GqhKENw8g
f3Mlha497KllO2I87jNo/ozU6NHFCWw6kylWSVY/T0rNe/DTtT2okSgwiRlR6Fig
PWaLBBu0WyB8D5VO+VUcWKVzaCh3HyZtIQM1oGeI8pxShBmOAKk4AqgQxdHVcgtZ
llUQOfsfwE79jgfCc+M2K0vB9OPBqHsNaoflg5fg4JGWCvipY2/rMrb/MW7nFe/G
Wap48mwXKgVmykgimrAixzCkUl3yr9xdtSWLjNVLVdKTgF7LkY8ImTMiypUVcUNU
7e0jCDUNmNTS8DW1Z8V/YGWm6dLDpcGylgus7pz+W48F+z09Old7PSOQCjet4r9g
uucQIbJB7xzBH4hvr/5xvWn/4/zAxnMbCdsATtJe00rQyMWX8+L+ht1pYESslOY7
yDbO5Mb+ZFa+VhTUda7cR7UWcRvwLxfWHv1Etdj350ifKuxiiA2nVHIQBStllg0L
lN4mm1ZeRBzSrD5uBL1VfiCr0EH6DtcWv+uh2i7lxbDjkDkAY6wOlsunIjr3pUGf
E5Bcvm7RnoXsxY6Cidvo6QI8hyo97p50mLQyyBSKE21I0Mi/AJjNHwNukPK/8v55
LgzWNLn2aI/wder5ukR3JWuLFVDV6wMqeDVc+++8/EA39d5CUzvpI5jcBUbOJv2k
l+VqhHFPcCVfZfxciMnJ6rmernAsl2zNYu/hLu6GwCEVNK6YE+Ofkr3d8SQxKrJ6
gaqz17UlcqyrUBqjUpBhhcETC5gOQ2C9xZbnMtVLHF+qjkGjW9QqWeTrXdxwbgeP
a1IfDuGposcBmoNaNB5uKt942SFCpV3ZiomZS/r3wqd0GhtfE/iP1J5dk+ck1PMn
zswkaK4RW6dfvP/v4r43RPH68/Esms5QqjVgQSOHzxxneIygeUSKxbTPLVxiGYDj
G8/32Qw4BLzPSp934hwVDecJS3BrSsnNibDUda0fwbNYh9DDDE6RWJosiwCY+tXY
fCQ8+97riQp4/KYcBxYNxcOgzeivDQ81k+RUB0GyQW+4P9uOgMuLmLuBT6QSis1V
AJEOC2ztGbRGNasz+Vv42DdHrsQg8NiNMSCgLYWkC7S7hgYtzfGkur52OetRsodK
NI3yKAODCAaj8vpm0zGwogwBuRwyOVkPCC57/FLnKr/akrUfqKWhljPDDCZ6hy8U
UrfSCDqDCPerkx4EAkZkSd3qD+xJ+yTa8T1xRPihvbJ0djVEpXjBO5cyqqF3Jp6V
aInQ7SvgbOtbAZPUXF8NRlD0kaerI0N2cixeLpaqobrDfC59ePRGmO/q2VEsLJKh
AI8QhQR/1aKeWngPixHfo9kN4olOfoOgO0ceBL9RLtw/A8a8pY6jfZjK0h1pgquF
McHDN7KXcUHFzzDVHld15ck/qyD2k/7Yt6/OaHJbbg4Wdkk0NEeIdXoXmIVYXA2D
2MqGLd7pYSPCGN2pF1683No7aIqOTBeH4yRozfVQFE11/UHoTG7ZhqkTl2y1G3bo
MCgsCQdikI2loanJyr76PPvSh1rFsnqSAXVJr5pfcG4Td1tfziMP7qZSZcTwzvPN
oD6XLqEojMLKHGzwxZ0ZRP/VOjSW98rWhdq5YRBgAz48mE+eThmw4IRPXcFHyvNo
zVclrmjc5r74ItE3aKSH3jqRF10apadW0g840WOaAm4C8hNOdR0x1ikgoJBdMSGV
38+zuBk4EWzpV3d8/BLBqE/ngHXe34I8lcSaItC6R1JNaTiXgdSNBT3l0MxKiBa6
ebqe0g3ZJByz4L9+zK1rl3hC3dCTXEgu4GybahzihgLdIgPcJT+GlxHgzJDq5t7x
JBBukR1lqj3YHWS2gzwvP4y1Sy5ki2OxVEQZCsULQ1JFOlE4poksvS0aok74aA2W
cgNLi8X48apWC6aH1A2N+pVFsetdadf7XjYH22ycz7HEx2ogBwxd3eroUBMo+svl
RwEYE0qzDy9Pd4JLd3pCgJFqRWOy59eTA4L9Wy5V35lg/GGY+uc2rFzBXEEGDZjv
EeISyy7nN6k7pRDNiSEEAd1hTSv15Oolk4e6mMPdHwvtiHIh9ZGlzFblDYms79bi
8LukuMsoebgcVezkY5b/hK3A6lyYVKosfCtI2zenmulqdFxHWtS0DYQ5FDBHH57f
lVbyqaMBRhhFvCZ2EWN1qAL1VhdQjGvgGlgLFOgTXf1jOZsDnsB0Tercf4paOZXp
4yFI3+U3ykwLPT6AQ9OefZnPmplb5N6Xd2ZO+YTFg/yL0knmuV+QdwIYBdJT03JQ
RPVaeZsmIM8PXcUPVppl76Abz7FZaV2rn3/QJbA+M/wbDJhbsX3QdvIYQYwQXfYx
Pd5qcumWK6eJ+KRV1/WPtOISut8W85Baos10UKufzvf1NRdFhH2eyGws/dynBrYn
IDN9+yQ1agFvIM9c3Y5df02u2rWZbHrCbWFHc9j9KrO8cVq6MbDwcA4zEuOvBeQT
QbP1OnaHIwYlmEOJiS9ITO1xIMxDFQQZlXDUvObxJI4CH/hNQGwSOzDWqP3qo85M
3gmRFhrdpUzVi+Ht/OivAkLDX+w/rgf2CSTrdB0xKgcYC0SDoeKvbAZhxisWWoPS
z1zMmd97U4+p9zG0qgcS7S2LtVYLjH2Ee/8cr9HHNICVCXN4xS2iQogMGc3w2t5u
AW+dqxDrvshLPtZv/h3N43gWYdclgJWTXj7VjuMwVIzfCpsobQ6wurRFYF63oEFx
P/hgLwBX+/btaapYPPTHNJrL3Bjo/ShnPeGEDTllFE2h5ut2C9Bk7sdGHolbRC1i
ch5AL7shO2uwCYK3xswXQQfIUUUkGrruidMSHxgt0Lhdhco51RoOICQMMYOFOROz
QAT5hzBM5fRF2sj9XwRVyvcDLkXhr51g3dUsFWOmEFGG339zEefFMs3q0mfNRrWi
mWFcMarHprYd7lcI5G/Ovw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Ky0pMD/3Y7x+Z9nrelvJ4Wn/Xn5YIuUoaSH/TaZJ3LfdHP1m8Mplf2wxRxnFumLF
p0DRQsc+eMabos5aZ+3bwIxKcYc2rVVBfaFr3gggxx1aGOWV9GhpOxifzuXo7D6b
g5oV/nhlrWIshORyTk436eCdki5fvf0XHKvkTyBAezY39PebR+7ArGdKvLYiZv/g
O9hdFxlpiJ7Vvi5TTmFN567tu53moiEqZ7Idz8XhgGGux4OnXXUUW0yougAhmsN3
fUjSB9naY33CULt83HuPmCGssSOb+GOg3ZSzQmhyzsauZ857s/4MVEI5n/hVJAwR
0UU3C2RnaK9hVN1MKNDYtg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2416 )
`pragma protect data_block
peADYMTzzqD2tVVX766oG0JbgpojhfEaPC4bOr0EwZ4SK5SGvNUYpVkHY/VgNf+z
T2WPw9spmQa43rARCSAQl/cSBQ79y8QbqyedQxDG1cPqk1Otb9e0eY9NVJbe9i5M
R3ynE84J3cDYnAImfPW7Vbzs8LqsOqEpztLa+EpTYawQNZlXSofK170aVAq0rHlX
zHj8gojB2UuU98I46SQl1mQ05km0Fp+0oRQ5NlDxHvt//XR5wNbPonVcxDJ5OZ8J
09u8zLHv5ZstOH8BYHYvNKfsZBNtraKIyLWzKzH37bb8c0PLxKwYt8uVw0gnwe9a
/XS485b3uhm8P55pn6z1Z/1TtR3EZvwCcv+FWcsmbHxo6UalGgy9XGf25D/wJa8I
98SByB/V9aEfTeYCRXCCnFCYpfXsm1rTWA4G2jzcIrfjHH8RXnoTJCWbx+GhZN24
k2jcNWTebvLW7a8vP85YLPMzyuuasOOzY0f0wAVvijv5YUfpAI4c9JD4psyz4n1B
YuIlTIAPFKMDDve3vjkFlI7atlPoWReR1b5GmjxEot1nq/brjoAySjAOlLAM7Wfy
SQnXMO6qVy3rJ+MIrogYvxiUq4D6p7qKsUkNDGrVPOZLMdRhterfRiZKkhEvP/dR
BouY053hRuk7B2pYp0LEoaO1Zbvi1ko0NgKzNU6p/m9VzeYslqz9an0dxCLxkCrN
Af0cVNJYokyoDB+Z0MhXJGlinlhFKkrUZ/JCR35QmcsXhop/AuAOSpmgvj3+eVmP
4Uz7ejfk+jMd9jmUsgfFPD0rOrhg1bTmj+yD9I7zXUyKzqkSv009M4qvbUV20lJj
0QbpvWXPcN8KN3Nq8RkNTcODRr6rAOJkxQo2nmFk7LRaYvQWZiMhj52HwjNYrSWG
VTiCQnJWF36KyuieVWBm8RETC436rSOt01C2LDosdpYoJGUo6wAeccefvKoPsnNP
fBTFO7dflbbCaLwcqR8+fP/02DnS8g1qqI6NsO+s3dfkBAXr6B24DdLiqU/s7U74
69xMAbP8l4Skl8BVYOLcN7WEumj4on9ziPEXraBBkZIpf+FyzhCM4Rc9pRiv6D+e
PLNhqrGD8OtXzENmmTIlqRqh+kqL07sXTAqZNkHhvz0iYRFz9sDvnG1wxlQLFw/x
vTp7l+08Dz29/mU0dtoNVHIRNiw/5AXs7Ma4TGBvULJZSaapZraLIpXDv4a80Q+d
/crKCIy3tDDSkPO43zfJ+tny1u5A60iLpgEHMwNPucDZisIGosUT+FrsF96PaDuN
kMa+GpmFTFPdPL+3EYvwAC3/jccQlrVVlXP9vupvpcHKFz2CGveRHbozzxSpGFzZ
NF1ElnbaAotiTonKvsu7+bcTnOikTyDjZEWZA7wYKpuFc9xy9E6VS4WS0YUc2Rvt
3mKhsaOuIXKAGvJg0vDxdH8v/DASPlRC/S/7gSEIwBJ5SV/b8uWIrDnhicmKnzmo
18eMJ7khkGBZcdNDxd6gXgJN61xjsLoSNKdqkRjUI+oNi0ciEDdo2J1/2zIkyxRb
sh9/wniM42X0oCFNEQv5FJ2GkGS5ga5CAdw9dY5Xt71OqGS4VXPfJcgWRaA3UQ9C
RcVxNd3+K0RwuN7I9KaJJzeMNA0ERYuaI0+ALKivmMvxV5MW/9AAyiYVpoFhkcE2
BJ5qQwjU/+uDdZf/ndSxoPu5jcsE+WWO8LjbA96oooOKoLGpaXA8zCOFxf57OWBa
AqEJp+jG355rhvxPloctimyvKXhUwZQPG0h/DEYeeYyvPuV8P5omnql6wESZdNDR
7kJ8Vd0VLtb18psMs8kvrHGpsIUILAs0OrK9tmkxyGrLp7OlMgLKxjOYZtWUsMRR
uaGjfBchthkl7sTZKoj/Treo+WWCodeO5rA3U19WOBmEhfUVDF1nzhgeJ5DFEcJR
wV5Ylqg4bYBPJ0dUSerqVdDvqWEyeudzwhyRgdHj9shsG8Hray80T2L/BSVo3oqW
SoYH2Dcdn15UucSl9/aePJodvXsH8w3gIYqnytIP2H43+Ioxbhewo8ZZ+oJYw/RQ
Jh76qo47UVVW6K1jGmcFCE9oWRnZZ3B+SekIXJlOx/SVDUi7XOZJk7wSvoUWCgSn
Hc+JUNbBVgTgRHUzobNqp5wopUFDlWGZMsqEPqGjQEEic0ISEsFshxDp7LOVXgpm
vkMGvKkNc3+RzjXqkeRbQIdR2gvOACVlIcLaxGX8wOKRneIit9Zw2viJczBK4TeH
UEiNvyjwyLW5fIsGxRRPg/UEW4/MPcZCd0QWsJEiDEQvDYcnip697rs6Lq17wSML
1za5XSV/8M8SZbXgBkWqzc3U6szL/zxyFykaTTtzNTc18fZ1sKqJ7lFlYujPTXmt
O7/n7FGn2YYuDHBvkb1m0MDNUrsDlCa8Uv4ykqx0Z70YgikNIoNAhm3+UGWVKM/1
XO8QrA+TKqh4jJzoo183TWKgRDT6w7raShrDlPXKFxWW+/8na7sRwvMuMYou3KiP
ECgnzdB71+uJCnzdl+tUSCroGcyqXMSlsfcxhnNYbjVrX8AHBUFWgMPM02WEYabE
058NIk7oy05yiBMlTV8+ba6GTbgIcN2QKMT68li40OQhOW260XqGPK7JSH+5y5qB
aLKPks+d++f22etYkdx6Wwc1hwx9D/R5ffHt4ANXajICVURoQ6o7lRrsN5Fw9dYJ
wSHrsYzLNUBbjGgwVwR3g+esyMmE4If9IfoXOKKt98XTCUiwpC3zi6Ai0o0xQaNx
95O8CmKN0PBms6t/9C+ZWX6r6XQt8j3YDz8KlPmmzEoWcWK91CK9ufkqnQqsCQ72
uGBfMmkR6aBk3PDoyld9k2LdD7y+ZKAzWap4p1VX1zDa+f9yCijKKGi7w8IpoaI8
eAlayofcfJo7m3cmt3ASFWmeLJ4+yxXBOJwZGgnIIArWS0+zlJxjEOrL9wVqCPMN
GrUr5Zqq+6ih51OFuwvTWD9VEPONqFmdJb4aHoCqTZctqpgQSGzK9cyFpElqqOgd
GU/gm4aVMokwpcAx/dpWwwrucIQ9AbCz8MG8CHS/kR3q0W2PWQ3ygi3AhRZIvEXk
9G+GJNnf9I271m3RHvq7JajlO+7hyOb0lh8HFA7FI8uEFA3TXyLwo/RAeL/rNMpp
Ps/du4OU9AUuWFO347PyP0s3ZKwK5DUshT2y0bodPD8lT5g8SJrnEajbLtBC5JxB
K8nZVuvkmn1t18n0Lt6SUQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
NWjRYcs+SqBXOpVDT98WlSe2D5n+A9NrQMbu/ZYVx7wzB2naBVlQ8lvThfi2lcXM
NGLPpVBP+BJSKHMEgw659ImqBC9O8bE43eHAEtcySpNrSlIJw8GsUk1LIp5fmND7
Fq3j5N6oNwvXKLnh0wKtYc31+UMFldhY8Eo3fjxlEmry5eYHQ9CVpOjUOXtoPkQq
pBLfI9TOOhLBVGOHDcQIPDhgH1kQW9qn+z/VCf6KNGR/WOqAc09fWpkB3LulFRWx
a/Y50mLD9N10rMUJBS0MWPH54l9k9hgu7UkLJW6jqvYJMIVGeh7DccYLBDWEjfIn
hPETRiokNjCRFZ4T84dfkg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1824 )
`pragma protect data_block
EC749D/FZHvtBDeV+0T31BrRFTRdmUJVti9bJZ8uOh+yo8sk/Jq2xdMV0V0SZnko
uFcfQamquLIAOEbcpvhotnBOgz+OcJyYq6y5zCxHrecWVuw0cS1CiToYdx9oy2Jd
9pba2WPVltFpY/K+21Oa9dcBJm9aLLz1xhh4SBKmf4+up7BCbmQbjx5ghrhKxMpo
bVg0ZmIpEc0RtArfWL2W+rC9eBlQ0bEkh94LQi/zTfQQw4ecnQA1Zp85vTpGKcAs
NKSiYUupfh0RlSORRaadfcBmjvBNy7A1Sj48/tpIBgTZDxKtOYGs8yAYDkyPGmZq
p5FHnk0wDDuUvF/d4AY2VBsFXjN1Y5UDkzPANITlhPDj8hLSUrcEd+t8Ib0eYFGw
4jX+7KYDhub3oZEOXkv85qtJF8W6D6pHJser9s+w95qLI8qBdX/tyYcTVY9EVNFL
ZibP4W7S0AEsHLxL3jsqlDlZ2M9n+92jfZ2AWxjMALRotB4t/amKsJ3UkSNU3V07
k8gTaVpXrNq5BDcHv4Sdo/mO1pvAnB/TdWCOwJe77HixBoxfoRDOzleKpnaEZDp/
KtyaUwsZMS8rHZ8RXYBKXLt/kf5WYezoBaDcbIcFCMYpFAzAbcnSmbfXc93gzs8v
ccg2rIBRETAt+pNrkj1w0HeZnof4hETH0Lx49R5y7PaZjKNL4kKL4fuQD64kysIu
MjJMgbVIe0DPbmSaOcgQp2bq88D3r4akYfl1VJ7kFQ+qk/9ihmKtLmYAUqiK+wKS
Wm58bBXfOMzG+CF9bZG7jiMTbGfvHoHikVZK+9epA1ePEdhmM7dG2KeZKJEyyJ+v
7t/vkmYXbdKDPMlIkwzYzMeOHa6mVAa7kebai9hRyn1ApTiCUUcHng8B+t86BuYh
GQAnbUDTNzRTnegdcH6/HEJXOO95Q6GLHYI41NHipurnC3fZR9vsvCE0CwoDV1zo
RvhdEnQ+vCEE6s+ckrKMxxjjV4BnprSAA5bdXpo0iMiR1pvTGviD46TAHlMobSUN
uiEkH9gEVvQWDGznaK4UZnn61WSSktZE38Z6QrapSxP+mEgRKySgZ5iBBTDdwgU6
h9PFb9+IZYJXMWBpKfXj4ZotWi/HPAc38qeJArZqxRfQJfV/Y9blqV9FbvojmAAm
JboMFz4j3t8CjMWJJg8A+Pm25h0wYrakBlHvJ0RgnmDL/GpzARCgDFf2RTHoi/HC
78IuykUrlmaOLHYuINCRVi3FI1dANceMlwoxxhtB2hvhrC3BhbzEqN5kp7D8GHJj
guQJEtJL6rRCz794GAGhocQONEQkJxrjqrFYAwiJsdcUvf2fTCv+v5HNdo/Efrms
w094nYHWE5A9hOKd1+s1LmPCJjeNZjUh2U7Cb49pYxXrcWNi6HM13n57IafEOxBC
Ql22EE2PFdoKhYCunGeKlX6F33z/g2gbS8+X3XfGFA/d9pvudOLOslFWMmi+sl3t
y2TzlxZ4k8qsASLXyW6DhaxunUcYsu5qDumjLmQ/QhPYT0o4Rigdf9v3eHtSJyuW
vXi3MWlWgfLdSBqriigYTlT+boiC8PVmyyx1Rgh5qAWbJhC+gqGj2j3kcyl+t4YR
3Y3o8gtbIxjdw3mOniODlTgdADM+tX2aeoC6Ts3NClwXNVYFXH0yu6J4jetYHz96
fP5qYnuPbv6YWQ0ryp5MfPlVasIEToX/+b+2FUooklD1Br9ef5H8qLuKEDNGadiD
fHyOSg4jyqPqBpEXYi/W/AOlVFV8a4Of8wAkA+pBh37CZ0PtDnejCAagHqXCi4jU
iK+Xv3soixPjEU+FVBOfUokD9pest5lfXnBE2tPqROQKh/l2g9dH+VLj1ZmjLFiL
wJyvG0SSnkFvaOEQsw+P0HhxJxMclmnt5syVudEkKzrKPgCviAtJvmFx/PU9Ke65
eTq0mzObzJKRD/R0+dyJfhvufPTl/nA3BFByovJaAvIdd19x4WFQxzUCquNOpOAL
2pBTsQguj23Fn1QVeFbt83PtJxVVI92AgFZsCaNrbSKSlSRPFdlF6G9b+HV0el6g
MKZmOeeTcDt0zOoSj0cfQvDl+cNX+hoCy7iU7xQKwCeNaOh2QmiXVc/PxMh6PHCA
q1bklygS4UWfmfqJdsB1od5XWWbG3P7d86UvqXM/wjJ9kngbb6SNfhCQoiInx7o7
u0hKIVnYr5VgEZ0+3b6UtBSiTMW8YI8YmmVkK7s/pcG4ogLJl//chX3JbvFecECg
CGwGW0CQwupJ206RSzSn8GvhAAeTw6A7Bn1BaUWR5/yzSs+53f+k6WUEEWPJ4c/r
xiZo0cM0y0H5EIjxFmHh0GbF6SLNDOldzoyUHGQl1NmSFMdZdmcPqhASMzFzthNy
Ap78dZ0WnKmuZ59PGvi4aah8wzndDGJjOVaebMQzFDKQuyTIZrmpRVJYykTIjmv8
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BVu2Zabju13dbU2haT12cDdXAPm6XQvqJH6Wj8WFQ62DZGG0tPdlxFPbjXpURiv8
DIKIj41kmzzWCxZk8Q1cElB2bx0HclnO71asv7ef3/LaVOfGXweHV9FsJTW0RLOd
M7ZukWQksXXmmn6y2McIToQ8HgxhIRSuABamQtxUJYWSER5q3CYyT9IA5kRfxxVg
EJtFn9GvIrebtIAx1sSIFFBwr3jk0TvDtnajqQdeWpu5a/pT92ekHUSZo3IbPtx3
JdqQxmXhERN633swy6B1pJ/QPmHm2oYb2ib73ACJCAxKnL+DsTBGisoIFNtx4v+B
7fm2l0a/UM2DTRQn++cgng==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 56416 )
`pragma protect data_block
2pZpM1APiX00p2pBPa3bWNFUhNrU4RqpwI39q2J/EWGpVSEDeUJVV680lZ9eJY/k
UGgGfQFggkEgZngDpWHGTCqM9g7Fo8BW5pI3/53LrVd5xiWURYgQGLe1QMIrixWc
G1QnHGDA6yVEZYFs6c2sBUodPBr5cqWLxzz0PuGOss9kx1O1xaT7p1F3n1/e40k5
9kSEzKdTLoSCEhaSiNTlNP/6dLLczy2UIf0xZjRLUpzmvlIsfenMnKeQoNufh81n
oGJ+YGZKQp6nHnUMj+UNL0gDbd2K/vVr5I4kOmBJolzw//psDna9wdsKecylWfxJ
Cs1/9lt2uD74G9ZsqhyScSwcwfTjNVkfHdBfP947aIzvr61LWGKChqETIX9J+BQM
1P/jlBF+6SpvFDVqqafsTNApiFCuxuty1hODIFm+9EO5jPDkGo17oEeYYYB3RlZ0
Cm/IKOQyd8Z6tjm9WKwvYo07wPkRBxW7sQTraAPp9uW2Zjyvdp3ujwUj0dEXf7dG
cF7TbfH2KgYR/Ydjt16oWpVEgoD8EnB6cwtx4YkUmVYRMuk+KgEMCl0TWZlunbZh
TfKPEZEnegdN3CJUmOmFNE//2vK0DHchFg1mbxjD43Yjsp+cy0/3Fe32P6riLGAt
OjQWqnlbEROeQcTHEta6mJEtRRrXYZHQjj13TUJjN+oMWqlkL8v/8fk5oxXdDfyv
sS5Yxx9iq2zgQlMJPZk/gI1hfb4ekBgAUO8HP5PZwE+XTJtOwuk1FijoXnYioI1w
afdPXBJutxpGD2kYTjMLHM8CaHcEpWur3RIOwZ9kKiZIj1RMSDjpURPuEIomnDQK
gOiuf69Gu4oD9WjKt6FCEEUHKLUbi8XfxgGH6smzILx14kVEL7qZ5Qa1oQqZgdoL
EkDow98ZB12VG1h5jx4G5xaDNPtjEw9+yIeCFQdOCX0dIKYMRBWfnYWBk65nQkwG
mOdZzUZj0G4rnPBMKoAj3/HqjXkKmix9hi+LHfw5CyQuuB+6ESPVJJLypu7BdLJ4
R6tTyb48N2Z8T8i3sJcT1FzdkNsAOcBOoDBAj0Ge4t77N1eK2CXOXrZnsipE35w+
OKGzHTn4mPCVOkhMXPMhvuSzIFKyrxDBnuEH8QFQn9IM4iP6BIBVAycv1kOJmBqB
uBU1GJjrRcVwN7DBsH9gnpAz2SmGUGzF+2/UharJbqU71T8M9n6ChoNyO5mQTbrn
LvsFi8rfUgvyBcVDE2goXqkbQYUDMhjKtEGxEv536JpVTZ0nUx20ziFJMN0PnV15
5e5Dc3mVGcLYsHckvBL+n4w5LQYUMHfaqeosMG7iJPiKrk9La+8WkCAq0SbWMCxk
B6LNuFq1oklDlHZ+7tKgh98+UXU+NWRQaeDyRJ+eORLwOe2e55RJg+B2JkR5P2QH
hLQT4gPYhN8psKN5Vo9d5LhPM5UI6zY2EQCV6tKh+1afdv8gbapibtI7iZv7FsNm
4X0Kxt6a+yTu7QcV+qA8AfFmOJ4bU48xc6bCxh/oQ8q79XDMzt1G5CUB6C/mTkXB
IZ5qM6ETMyqfoT6cGiwAnDw85CDkkiR/eIfGSer4xk1OYINjy0lDZNzdtPnnMfkd
EaS3UxRk4JAsTUc5sHD6+tewAisZMPS1zIM8K2HiPietQrGFscEaJXN9zSXgOwic
NSqAThvnwbJr6Lq5u0gdFrr9j0JitZiCdCIh5rhesaK6hEahuIV9+aYuwPSceLnN
RvtYNld+csZ/tmvsnRORhvio2s33yZCG26G8g+LjLFdumi0nvr8nI2hgKabUyaiE
ES5yyszcRzwCdjwhZyusE8eoKXauMrJlMJWWcYtNb6/0MpDhV0m8mkgTPvW1Adoy
CtEl4wtWXg7ttwxKXkA7MLAFzzv1ivqQUaEkc1shKrasdzyQwQhnV/zvhUqdJCda
EsoDmULzH+1YypyQi7eOJ43f7VEy/W/5z9zrVXVQtjuZt0Z3qBPDpwHKWy9Fvpph
GJyQbeh1NI2V8dXg4ZLKCCIsD5lEdk4YfVseAwWAwayZGCMNV8p25BbYChBargjU
LMWqwnEdghLGCq/J28W7b6+SK7XpVqnO4oNJTsyFOzh2l9JQeViTnF5mDHmVzj13
mzNO9/1/b9u9sS8hDes1BzBMm3QEgVNThFTVfsxiDkU5L9WaqoZCW1BJN8WzgdQq
1Wqv+neUKjjycejnyOkiIMYeZEzjeWrPCn8B3+MZRasPzAPCUPCliUDBx1krMjdC
HCP+voPmDVgmm/ODwHzIuJPT64dZA71sIrMT0JfJCpjvw/z8zNj2d5S2Rdod+Dj5
UIg3FvWrJzor4FrsvH/zyGobTyvRlTQf/xQm7psr/n7d/aaORfo86J+oi0/+3aqo
Kfwpni/sdG3JxKE7EfyIqsfM4IThfHia+AK71Xl6a7F28fx1ANdeL01MeeK96LfG
G4imiAiKl+56MoWTr0GULuKyblGzBHjRmWeJk+ttKZVW+UDJ8xVYeKp/Gp4PflhX
zHsKjChbSxUsAwQJdbXEllf/2GPbGhgpGZL4NNmCWOd0zb0nN+b6nTxm8QTctKtT
VauZfHkASXkUzL+zye40WuQAZiRxzW6wyhpEFJGA8KuoddhmUGi5cGmcypprCL3d
QqLwTs0ZJ3VTM3OacVLADYXDfG9bOD/FhogMcxM/d20YyNeDu6JPI/fmNiP7ZpyA
xubt7kwStKCMMUb047jZst55sRw202TNqI3PdNzXkkXTHL7N/JhHpqgZ+jLt1IWp
epcR7t7U7bB+kd3mjO2FoXs5QUFHkUIJ2FpVGSSq+zgB7I45WQVU1XxnbZaFIV7Y
YHvuuCx7j8cnmvuTw4ah0A3+g9CpTQ0ZcqsItpwe0WDBTyIUC/gJhxKWQXAvOZsq
VNpkLnxrjWAMKOjCa5oLyHJJeVeYt/VkLrEXxQY6HoXdVAbGXx8Fllk9KYdNJsRQ
BltqfmTbtfwT2YAGbYL+TIYz/XxUKl4Uw7dRvsDXLnyAiP/w5JR7gPDBp5CRltZD
mWn24y/PvFNdIm3rZgBSwMKJF0llUwolh5Pt/GsKKGw4uIe9xrQBmwtpBjpX7RMo
YHiPwvAfbKf40yZL8LKW86GuSHCKqHmKt+WPq852sWelKZmk1SF3cbQkC+xewuaP
WS0Hog5ezsLNEDSEMpzrcnFKrzWJhYYN6gcjQVuAME9K24s2U+TqtUclzO4Z2AyW
snA6sBmfJXQlPqSP0xCDyikDD6SD2CaZ3ts0DympzrPFGDUcJNCmEq8fUbFBEtCK
5NvkUuIp0y47b+TzJcC6BTgFlSINxw8sZpeeR9gs56vCtXFWqTrINiAC65TsUfpT
hzsZoU81zG+xZiBSCIrpMdYtonK+RaexseIiIDG3H8eh54LqS9mxOdKb+wak3fW8
kutoDc/b/SXeeU9bjBxKZ4saaqoW1YNHUl4TsAuO3n2wwsBhDfrVxnwJNF/wUv5Q
U8z7GTDyPzOtSmE6eVgk5+chiJzcGLQIalw/uaCLhXt9Oxf6H9liVliJCMl9kjBU
PV4jwqo/ajItk4EVVGfBJLd4GM8mzth7V5VqHbkNfTvp2UleREnlUDie/Mry2bEX
ph8Q6eWgXGlASO7dACK5FFoxCflqYS4UnsXeE0wJbtBHkNrJYvRGmwqE6hvFbA49
bM7wFt8WEQzytcj/p3Y/UqSigncPRAyRCj5yNvCLYnT0p8osOmDyBwGOijCpK303
zE0JPCt8nE006yoEUyWcJ97Jhx4mdTmlwq4V35AfCoIFVvm+B+g+wDOLUdMjDCmy
smN+qcbDlQQP53c3TQx6njbggQIO5VxLBAzwTEaAlh5CJtnKpMlT8KZGthMxGA+N
JneZ1XNg5ccn9HZbOmDXzoojlQr1rNfCVAeMMFW2sludalfXrhhqOkQTZio+UTds
0BeS5Yrmpk5dT2lqWe3saER4DEpfEY4CPRXJ9AT87TOi1cmD3xcTlGudOfHIwlBe
MFSp+mFG9jrTDdpY0EFUXf8oyxhsniSCqb16ioAQ1GhnX4N9d98jMjJdV9nUtlq/
pflx/iJR7jR2KLsvd/6kZIPfoFQo6bPZGtYJ3q6Uy9smu24Bcz+ek9n89itrN2Bs
B4ocIAHqwPhgEQU6EQ0Dgnzp459eY75G0QowSzV6on/y9/KKTV9FVo3qG5zhHoJK
2wrI0PRqUAHsBJEva9fjJrm0qVOVVHr18jnhnDI9VFn4dpIbxsUp0vENbUuAIEC7
2YCCCn+azWuXNtABG1M1sBls2ql9cocN444R+dpKUtMVrkuG3mBhkDXaI7Klv4G1
cyhkd7RYWni9RlcryktIap9tX2mVhaIdsQFVJBYFi82i4Pu+Xna+ezo4LR0k9aC0
fdArjBV7iTAWJin8i0cXjgipevIWwCfc70syZForgH+KpHwusT5yNj5xWQgct+2L
7afPoKNTCe2/OrylL458rtQxyEETtV6yAk7wXz9UdljwOPgXE7XQRHXLsKq65tw2
WeRlpq9OTyI2ZdadhqqN9hpGJixJiqobLBZME+bGhs2kyeDdaWLIAbwkQEIDj5Ek
lyv4rSwxMMzdtxYN4+kNu/9frje9Z/nN3GOaDyY9+1/kR2Mif2Z86+PJ9147yuUI
CkWM/zDxY5ePeUa4fyzWMvP9YovbiPxreqgnGQfPZgTuDsEeh8ST6gMSTlmQUxQu
JlVlilsSwJg7mNXAGgsiAdpjJ2ryYx4z3mrlZGj2PQstI5xq9rERx/jtTyJkvt7u
nqCiGbm09rlQfK8nndIWcdT+XgF12XFFQWqYOdIyPhcLht3QyF5EK+VCfcqa3r0x
OXRHXq0ZlltV5rIm5Pk8HA10uy4sEnCyaR6EyRorJe24csIFhemFks40q3I+iszY
G63j7Rs9hDBwPg9LZb4xSznekBVKatazW1RFOlETiGW5Zj5/WEj02Kj6S31fStET
0B5+oXbcG0bMUYrW+gSEX8K+iwiCaguUjAZP/y8IzJsUCvMrIjYygBfpl1RBX7pc
8xiWY0UYgh3u2jZeCkt2xewppTMHmDoyfj92h7A/W3fpc0WrkwVImh4TZXCj9Nsd
S1ouOmyfJk2jMaX9Wh0W6XOWE9V4DyNmyijbRncjeg2YilzoNwWuleQ/Q/tvDF/o
oqG6eXACfxBHs9IEFXJcrrh5oO3A0UnqkHYbzF2cJAsLmwm54MFl1Ld4kG0Pr2bW
U+xiId+455NJC6+CGxDQCyvXQiragQuhI1YkzMVVA4cd1+XJrIY/Q1tD3C38DEji
pxX0m9kEKX4Luo4yz/P9JESXwFNur15a1g7pi6LdpMIWBI4Y197Ag+R56OdCtA+d
msyMD9/5KwxgyCVQuxtPN7FhxuLDJEo7Y7cJpOAZuXN7olizwooKICHneIGEcJp3
/VdmWLRGUyp6WbPCldTkG5/CTRgrDNq2bgeKjtkAQRWcB5SKuAOeNJMTGVCgSSbi
aqHRGYcwQ9grKNSJBW8o20GwwUut6irUJht1ppj4SBrtTQiYg4ErgOass+eFBvFN
inEExCY59rSYrsdUY3PSa/yuTdBmmJeRIWFsetckDXXsKs2AauR8URjEj3lLo+Qs
3zgu4sYNgx2CJRSgl/s09of2wJT2/uO/rkGE80QAEkVVO8Qr4x6sUmpq0DDXILoG
0UQzGUzf5vICVDMLos3XIfFkbHAzPJf5SoUEBXCoG8GmGOLhtP7ySo4azMK/W+M2
aw4q9uazmFC0fyeYD9UYRknIuTmXmfb1TUsbkUWuWmgvgdAe4N6O0Y1JeIVEf/BA
5v/u/r5YaiHm2dVLZ/Y8zD3l7jLHYa2xImPHsCr8Oa+M0aJ7Zu8iIb7QK14sNVaX
GbfLgmMjoz0o+RF4+KL6a8Bmxsg5t0ZX3OKYsrbmF6THoUi7G16f2l3U872Ibs6c
/R7AYA18tMP7rHw31zH5WV4dAhP28EHd/TTwx8xhuier3+nXBgrCDrlXpp0f9lnL
fG8aR4hsnmhG+MU/b9bbvF2+uKnR9nPoH73Fd5Nt7U6ly5+7WXd0cKdogmIXzJdT
cf0ixRo6NCaIiZRhC0XXDi7QLcXmxX2ntQ9/8pzMa8ChsH8K7fxdbhZWGSNU4Bsi
X5TecgTPBp4PKzx2gjAybe/xTc+TPx3WtqAB4r5Sr79WEr6NBaUOSAZbHwYCXVHO
uL+nHzDKDaMzved0ddKSfwI5kSbpPo8UbUA6QVvT0iGRMsJa3ju+VfEumEvUbPcL
s9Ww56a41kXF8E3kFV+vw4VbxIBlUIoqUIZ7pvZzfwOUyP+LyVj2RaCywMV1fIJq
MoKULYJE3WGqCJ+yN9mKU6Kox0ysW3UHAQwzBlFP6oA/ofhfkrV0pFMbeAZXmAka
k7xK3XZpCFUxy5SZ6pDCKuIE8SvIkwkQuKuYhxJ/jfkZYVUPrv+5CbwU6m4xPq20
WBMjqEC1BQZwP7YLOD2xq/FMJknSkCKSs2eOWTgWP3Ahp5eYhaG+d0Ob5zELWHt4
+oSCgae/L8R8sc5CdxgFQB7v/79RPV3IZ0KunOxcYGKAHmYtRCOCm7Nf2pdozfwz
dcYMs9bsXeyEhQCnLQyTlllh4KIXHhFKAJYVy+8YrzX3dYw8SVjjNM21L7Z9aMro
hPAXzPP04L57A5YO+/p7guTa1yXJYxATECnmh3rcvEqYAPeKE5bfOmb92R4JiBBr
U+rEK5LBdOMpUwsh2iNezbHfWLQJqF8U5XGxddvQGKrAiDKzUU9ffPyZiYUCS88T
x+w5REiBz6gUXL6dqPQUwEPAD/Xq/sFTNuCNXOFZ9BIgIXmyUdSorShAwmCt//Ly
RxVUKLUDuP7+olvek4xMKxVMgKKFavdauy9ovJ3IRkCovbEblztLo0+K/Cyf6eCh
SIw4SDYLWjBWfo/3xObXVRguToCpFMVVvAzRj2UoR8RD7VpyeJ/RKgEbT88eOIFI
pLUlFYosMrkXUpzyDRvqalktLKxh+PvnSgASAvmrqQHPsyJLvC05FBit+RlbwUSX
R9Dcy7UHymMmqub3Ur3NxvpwNIOlkklTLTivLzVMjyM3N+rUX7T2OfvE4NG6STQF
QYUfGUsZCjc/PIMe1M5qdIm6hthdGYkgOBoR/o6t0DUuTHFyKd+6qxkW8UhUAunQ
462fmhivxrNma7Fwq0PIKI1RDzR/He5JLZeajBFLd1H6OV5qXMWZCWrMs0PTOme4
ofAch5xqlj9AASLIzRL+3LHujlbCj+n9S9JtDORGI60Rk/19kuCjh+9qxizvD+db
QjWwXmvTlq9C2lmBy5jmjSk89H4cwfCv/lLBP0z9DXi4SayLkVQrwEzdjpv40PQt
pIGd26IZ00I+6eCIySeHSs4p7H5ljjY+YS+DjVmcHx/SZUWHWAPbhFiBKuon55g0
f1zgMqLRHj9XUK0G8LVGGkJic0h7mZNzXGV7wh0xLs3OvS7ye9lq9Zerg/kUJXxm
oQ8ideT98r5OYu2TZikAoZ/ntWsKmWqoToR8TzD+uuoWyCnsC04YzgPzi2xz314W
8AW0dezl9TC84DOdcpHfDmB15dS1mBQKarbEqHN8/e3hZK4V8/GgQP8Cm74NiTSx
FIXFZUIiDUaQbUqgyRgtlka2crM5EYKkP1CscRtVg9Wq+DkrcNieUruG1/bsyK0K
0AfTvxxsvgCwWYNBu3Fed4nBuq9PmfyJ0vR5tpp0oC1k2wuaTqpd0M+KT/7/TX7b
ZSMIOUWjbA8p+5Ko7kKd3/p3IDCqsFbtc0N94clKD7w7AXo7xLjflz3yVXiWTQCp
DT9nwFDBah+8m5P7d5/jLRDlvn6FrN98W0J4X08SkNwlmIQVLBmlY0xxdvYeKzAH
FTttkTtnmzTGDkdVyNPNVrwk+6OHhMaI4QVs18h0tl0jSA/9QKOssGsZV2Bu278U
baXAxXKgUddffHrRo3jq4D0HFibPNiimpJL8fjBwI0JOAKoG7vXF2K09CK1c/6Bl
zebBIFD6X2QWm3LSr2SPfUdEZ4CrjIbZoOxxEpR8vJMUoxNdARW2LbeeKqZrbl/6
FEd4+O3OBJqkzFV2t5uYyV2IOap+kgZ+GuiLa+hkpKWOkNE9AoWccfaSoxR07zFZ
8Ox1exMZx57XRzz4Xz6THJ7A7JriXuLGXM2psK7sAGHACvTvPh7EZoOlT83mKb2a
y0yOshgMz7vuResl4iOmTb7SyKe/4xxw1CNb1OqBo/VVUntTyUgl5esjY+isBBIy
0wr8r8ZTBfndS/dsABc7kobBNV+bCYdSJW2+m2VYDSvj+b27cM9SBCFj9JixLUq7
IN6r5ZYNaGYbPnqqeKAlSXVwKu0mX5c+ZMNL8TLRvL0ly2YkZ37bk5cCuAwbU9ZQ
1Hbg8B3dJCPohLmJiXY3K76eWSARjrMgcSiHYybN45aMM6b9xaCXhTHrlG9it3pl
uMRCPsP4w0iSTesaiRgLa7a0K6bwRov5KEJgcr2XB8huv2sbgb/FI5jojNVB9K07
T1K3aBDjYgrW88JiBpkwgjJ4mdkVJ7p5XDvgr3FHaHrADcg+kKStWqOrUPuN+Hn0
z68t7bhu9JU/Ng9+nm/s8C9pXGIBjHHn8N1+/g4p0Oe0VlDDoxxvM3adY/1pi9hi
uIcB5vPegyb7VDhUaqsZNpNruUu4x4wubuWAs5ziPiatGvT8u43BA4n/Nn9oSsYv
pjkGOao+sgjPZPzIEqB1DCHb7IF/bD7mgfIKU4AoZLj36Fib/KnkJFtj9wOFic+Z
D2Rd1NlNrr29DqAQsokpoz8Q27KpDYJ0KjG80B27SswgMR86dS1N7vIbcrSSTFoP
QXiGyRVh20A8tEdrJnpUYYQujMFqbJnfNdbWDuaYICD11miTl8PiP/oRDu2pPkhH
6GeDXq6jhiJVPZdgV+qZvWoGRSz7WtcF3btKE25FmmgQRwB6M7XCfCYnnFmXo3ZX
k0qA6nBlddFF536lqt8QMMHEgRlJVVFzASDQNlu6NZ4ddM3oa1vVkkzX1w+G6suc
uEU6HWoRXsGcWP0SHwdeoihbAtRv1oGuVRd3J04oQbdaP0Ah75GIXJiyRB6yVT7t
stLKOvvnqrS1vzVxLvsNNHQktvpRHpunpVAsKTjIxeuCVkj1Tmv0LnNjbNzMGcKP
Z59uCR6YIEFbo7InL9YCFJEBgbfJ5hXc85irU57xBJd+JHln6g6fLGOf/XxTX9TE
lCC9J6vXQ/aZmHJtdCqBGD6NSPeVnIodb7e85WwNCk9lmlgPACA5elCLKie5F61S
98EOEvMqU+Tm3dEsnzOBwdYfAklmHw+TeAoff1yZmd2Xq1Zh5V6Fzy/xw3hcRK/p
a/zTAYlggnnfqiFMQ3oikqkY1kBQsyJt98d6cqK2DD12QM25aPZCC/ZMnkRtqkuV
Dk/kfs4nzBP9OIjSy8JduxTEMTqDO+go0KnALxLSSEkP0apuHmq8nvq388gmsk9V
6mxpGjQw9yMBt0eWoJJz1K6gQSndLKfiCtGBLX2sFzpSbubr9ziYuyMT8BgHwHQf
jSpvEWjTWBlDliH1lbXMhYWYWYUh4L5eg1kobtFck2MTg3JuTeR3n+Oi+lXwhCLc
pvTUi8E6TULfZq6JqLWQGLbnrVvBdeWumCH+ile/U81UsV6EuU1m1+5FYY8HbTTz
uEAbHaBWaIEnhI4UHM/2eDfebEGTZJCOtjyLkCZsoYBw4thwjYNece7UcvD9NL86
BNgz7vNgb0SW6gGtevs+1Al4Ax4GAl9+NUcou4uTckNoKgwff8VDAlxbQmF4YurK
4X9m4RlNOXuuiXXtACAJToC0EO6sidqw2qFKdoEDfyRCceRL2k12W8njgd/oQDVW
KZfNTpMIyDhtEdZouEqC+OjbiwkKqeih0q46Kc40CBAod2yYi26AZwQKGG/uQGwe
J65S6s4x47+r5yZQQGZLYB54Lf3KqbYIoHlJ4B73fkdZ+IqWH6u31RyglBZoyhOa
a1IweWbuNcX/nGRKzyb6MxeAB3sngooMs8J7gtSVHLFWUoz/zxSPXNTXftfR4wH4
mYRwp6a2IFw7UzXGg1Mirop2JEBKBPVIUrnt28SmEKaovcSstHsTERxXnnF3wzEp
YYI/PjI8u0v6hpXRse2BmyjD8QqKBmzUhQ9aoG4FyHRTSDA7CebJewkFWxVkay5v
pUg9auB/uY0ayO7R2CtslwMBJQBCQKL27ZOf8qJrewCHUPKMuGnXgNgyl3YPwgwE
6c8SZZxrq9hLHCCAhjUP5IWOZ08i2/iHvgshPYo+CKpUe7Gkw6M/yL5Y69JlE8uW
ga1xGIgHTtXbOf2YAbG9givOjqQhMNDKwjMJMIcnBPEtDxu3ZohVXRwYDDDh683Q
fUTLisKtOXnhrRl37pA6oJR4qNgrJFa50BytCMLm3JHMPxCzZE8VDgFkmorMiukq
wrXdQreXoauvCbz6kl9NoEHh5vT8sJ27Lfa4o+z6Y0oalCeM8HmJToYUPkBPcHG+
eZRqYhFhpWKQmu4PGAA1dtC7/vT8D5ehNwpChDQDXpK2QvwGaxCV9DX5NLKOlPlR
yP0J+sfPqLndNkxs/vBXvNYYWNWVJO5SdHpIfQxhMb4rYfKsDZuCw0w8lnFXgcWu
j7ZDGd5NIi7GTvS20j1BDAlieDEn7Ey0QBFB+ntL5CUAA3gUfreeMSdnwEItXuNe
CgKA1l31hXMP0zyOAf7SQSfKLxGkTQ/CCTaJiB1CAd2cgtjyj2n1Vi6LidRZVeqx
3HzkkUXDJcMl8bgRpTdoQjLwwQf3D0ZGn8h1e4XzL8+4htsm2Bjb+M19xXB5Hjv+
2Hq0iVvOV5dc3LL8ohyd/YzlQQlrMbVV7yGWfzkmLH30s7LAIT99yNIa9D7iIj78
ipOhxAnY5Fsqt12irWzs2KwDbAVAt7Xx3ldP8L8BTKlkw8DwTNX0hYpNVl1TZLx1
s5LtBbpqCFwwcMzWGqsx0JSIZI7jjI7j2cAQZplPJUQGorBOKRPXCs2uMPpzijQm
ia0qgpbOctqswR90nwCcmxbqCSqPp7fVfhbq5BPWWMXl51FEpvq7lkNAgwYiQFKU
LLNUcPUZs+Y3UVjV3ha5OajOBG3/I2TWe+PyPNHo3HYP8dnbbQmDhzlOFeb8X8xI
f0H9nkCx7rEVFRoFdMAaoTFUNu27hpMCwbEoQGZOjbjlGLHDEm2cmpJe8P9QdGg1
kALmcjhlg4V7uc8mb07L9zB9Ro0X2BTk5ZKq+r2f7y0La5hSeUjwOfC81wdKqJtg
chbPUtiFMPtfUT7es3fUETgPc3MPxQtor4o7vZwhJr1ceUYUgF84IXmTch8dGbmS
o5btMvvYGKdWj0pI74mJqrXuuuW9OhzVUAGoA+Ulj/stqwnBUZ62yVseiwvKIe3Q
DjwWpFJjMXkDi+ahI+Qhgo5tk+4dKHD8sIuOmQUpHJx3YLZ28VSnBUVXOXDO1KFZ
1tnZbo47umG9NmXlfL2PcxIaUyaw3xys8QX8rWZc6ax0I6W3v836wh3stTkK4k73
9toGJW+6oBQCReaIuO/x05TTmDgBAjAcDx903bizIciV9T7QRD6gRW1Pcpvm80zv
GX2yy8+tIO8vCxdXkkdLdwsUrpB0/FADV53j9cK+gaD5B2P5U4x+/wVTB+qoyxRK
Ur9iJzaDsgADs76oNPuEdr7mLOkCWp2ffyw7dC0f7+gu0rUm8Qp4Ct7M3qPS8wre
oDBsUiwKHqybiLIAKeiBmFWf8ftgBh3M/DVXoDlnqTrZMfrE+15tePP32TmDCQAi
NCcmygEVf+E5DxzK5obVfy9trCjMfqT7CMht5wxGWqLwInn7oHsm7JJ7OF1Ofmu9
uIhEkmOKHUzy4lAk4AqGImQFUb8AUVNivtbHmgmEtLXa6eTV2u/wl/dk5Tfg5zk2
LIj1ZKzitPblfM8fk/bRH3av0kTD+F5Rdgkx6gepMiqnU2HG34NYI1ksaFin9mPa
KUwk/zhGXIxhuMPce242sipLYQEeoRPElgnDmb6QZu4H5LMaMPvjezVM8GxIeQhn
0wEp9JO1tuIAIGNDiecdWwj9T10szFB1Z8pAyeQt2KfOR6I2BWKXGUsuTESrYtUi
5+xjRWWTmRrgF9LbcsmyX2snhcli0J/zgqWBeM7lbMLFixwtIg2yXGTdG91gYaz0
BRwhHyjCc+zZmvTiPzYYC/TLfAICGE3AX0CJFob9nFigzyxXG5eJUxPC8S/jgKXU
DIGgkE5AWz+w0ESxmHTD9XFhszf34sm1ElFZaZpJV4GpzWVTqCuyO4FscBy5gzdE
j6mDDPjJOCGrUPUxBnsN/4jptUBTUOEpmeZdrVhCK4oQsdYn4oZHlqCy3xb09qt4
ID0DqTziOqn4FwPYkIOac//TLIknZ4j2YQpLwwVQFEBYWXxmEsALYoZ3oyC2xFTa
Z3UuLvmcKZObstTbby7m6OxM1ODzY0gfdb2Cfb6KSOFnAB1i9N2+sVZL6KAWnSl0
GK4IeiN7yWU0gD7wIcn0203kEJR3V6CMZPN+bizUE3jxEdZtW8hbffjZzQ6iTPIt
pB4ydds8ZqDyPhjEHmHDf5cq0U34eFL4RJ7zFGICl/DyLl75e7aZh8N48jxc/EVU
94/oySB0Mr4jVPST34yhRVVk3QVG+1cPRQiCIcx80GzyORK6/g3wwP5YQLkDRVOr
oHHS+9eqSgOxLGj0x8ry+MciDWPxN5cwCj35JL/K/C419UeO0gFnVz6ZRg0az43K
Kn6lGLJ3vKakrKzvUfsLAl2SuS4sxUFE/GO7uyS3qFELBBZTVil1uGKICe9UH9Lk
5UtLicJx0nvGxez4QbKmvLxohnmjFTn0lhEuizjmL87HxXSxttXeldjyqRbi3TTW
hdC1wvYKSSUt9NCQIJOsoWo39MUx790Pps14OomCT/gFG5zlBAPyXVZukkY8hTcN
muhYeLdCTNVi3OYgjcJ5KipoyPq4+vFyu2b0Hk40lQz3UMD7BmWF2wKZbip2oUGg
d5i1zlNpKOFzdDTHHpXxQ6KVe+L3XTj93/xONF2iHpi6HWnpnhSj8SEQUrxHoVoz
+SWV9KunrgYFrYDJNWQWeiR2EBN09kGlVe6/SLBvw3moR6gRyPvcF5vF6HVIMBr+
GXC6WpYm2u8vcJVZ5gxKoCa9KzARWhA/AvvCyd6ophlwEXjXV+Ag9nW015Kq1VBu
9IUdHYWyvYxt9K5Ubwg9F+52cEPP4q6J8l7RuHm3PpCBu+OcEjGhWFlT/MXFHXlh
A9WewCX3iEf8XbEUeFihPKmsCXRdyLIfd+/yGKuMLebbbnTgW2TrV05S7PZ/rRbN
247VxXT1ZKGi30P6WJAI8xTzUfo7I36pwYSnbibK6L1lsveNRh0J8S0PGJ+4J37Y
1CyitET/W4Xslz56cXszO9DZK4A12+JsRN3OvB7Ysp+iYUjdN2WsefFrvBal4S1c
68XFTYqLfZZ3aVQfXk6V4csvpkE38bT9TsOzK9ky0q0wRCQ9B4i9DQ7O+Z99AQyg
CFaD2n1i0i6StTsqNcie2gw4IbtE0KarTMfqUeNLBfWB8ZXbAqa/NmMaSoZxjIag
k7MgqVqGC1wrMahisu/NgmBQeHtGrqEBZpP3SqlT9S7Qbmg6GcZZNhKqW/rFyRaJ
d+2BV9xqhI4U11OAhsjaD/+RYW9ZzSxUl2FHSZFsbv2pgjP6bkQYEXLZOSPKyYvT
CTJp6Dw2lHH5iavlDmbzSrkQ057hFmGh26IALLH+Aemf2Wgl/RcF+keHOb23pXIb
Pl1gsrFtpsd7UKys2WQV5Q8PJA/GTOwcwkUkJOjVNc6YWOEgTQkKBz3DSdu5Cq0v
35u//CTQnwfvh9Yz9bkXOXhJ3cAPJcb5SuRYSh3gxiYnU1FN6ZFrVNU3NwGPPdlF
uzl08w3KQf1Ur2mNGZ2B2rv42MIAQpdsLMrmL6pejGQNCaVzmw79l6UHjt+cbaBn
JZDz+3M3eEuHTBKhWfjG7unWDs+64BtGHc7Em5ZlDkPTnwgefyDDBE2lAOH3NuqN
1WvN3+lkFejvnZ99PHX+QaHut4I8THZEslbKS1wCr96c2eZcfEFohSP1sPrXlX2f
rEB1G1pdl4XjQevzi47mqJbGbjRLrzgpYimTA1Yj+EnyL/D7+RTbPfHGckfwBb1E
h6Jwi7Ovc6+XRc0p8lG7xwJX5Z5Z5vm7hBFYvsDV6fSw2rXBghGFjPY4Ke5qONWp
JZGd7pnlNCzFcHBwPLmgi6AmlFMJ3iaaPf3XFBRVLx59wsmX2EFi2PXBMq0DDOtc
jjA4/K0GrCVDFLH6WFHCXy4rkSYgZwJnnBapcfmPJRjCVXlZSYoNKYgLRJvfvlrc
Fklvh/ojp5yI1Q0xYXtpWDF4dkmgegg5+D0qidS/L/HCd1yn3+VxHNI9DNO4GvXP
wGdUx60dBrbvjxbtaLJcymZtGjOkJHRYEMAJJNDa3Q8+LyGJB+wu/TCYFLE+Nnv3
wwi7Pf9htUpyeXD+wK3GKLngF37TzqbYUdYzXf+4D3qOMqTrl8vVzgku/xB/Hf7Q
mHkizHVCXb82lMZ2ftw1FYg9k8HTDE93uJc4nPN8X+GL/ERtRMx7iQSyup6EHLgN
b4VK8fb5EIsrHokIY5nqvqMrVzrWxA18MqBa4ZCDHcm/+B1TrPqeO3FpDcj+cZXd
u1cjVtGFZI0726MG9OkLbU6Gron7noxDJ1jrG0lrvCR45z9vRbzoLEfeG3u4Hsfm
nikW9vfTbR02f1QjgA41hWj+4d7pBXaTRE6kSqrNP2OeCMztRaxza9go4Xmu1HPM
Q+xu8MfEAJOs5XyXbtcdTnPpD3M+ooTVQRHN+so15Ilhu4+M10KZjTPyKKcKUnA7
TrNhezu2xgBW5ui6NpuAEAvmL1m5zYrtm6fFLScH9XZ98DrSl2T46As4/PRHiL9t
SOroZcMeqD4wklwofaoJeWuljreEerYgjeSpJ0Yypthf1B0q+9cVtaScSek3nVlk
XQlrjccWOhV3M63YettqEE6rh8yEa+4FuYDILNwkSQKnoh1P+Qzs/rht3Rhw1hhe
xUZcpsf7xz+hBBOGGgkMDEKj83C8EBCyNTFQ1N+IfZ+sUfyLw6LoH/UV/Mkrc14C
Q4wEO2ZRXjVPeief/uGPx/2KZdh4qV+ftyZJtbBbbi0cqzlUXeVZEq3sloZ8lTYv
WvegCXAxpvz4e4qalq5dZu4tDugvuvLTEs+lWRQSYCNZcLEH7EYZ+fGNnb6XQ6Zc
Q+UBHlryhsjfp7W3EjNPq+tgQr19sG+9culxtGl6s9Lrlt/L9WL5BfGs43uotPXK
SAPzQJjtNlLm86/U5BkM7V1GH4x4tgxzUsfPDl+1D3o/chHHP8W3h0KVA4xHmTtg
ZjXWTcjh0cFOZ8eLv8VZXIiyKvqn4xOskBC4+Re8jT+9sVZ9bEtzeGxflv5ZlCOQ
92Xnz6RSD5m1cG+Q+60XN3J1cqDUPPYttU+kSmCYHMYgwaCUTg3emKLh4G+ASlTo
7Fzfqcnumje2aVD3Q0ye7vyih7DwSn0y/Mh4wcTzlvFBQ0OHS3yg6tEFyIQND+35
JViLqAzzPgtbP94MOHXbJeJ3L+ouKa36F2gOBHx/1tgMD0FmfSrUa1vEnm6J4G1X
UMkr1loCWKr7lZ3E5P0z9n0biHqVgLt8bPi+IzHc7BNXOtNIRw3kn0+bOCGLBqMg
Tp1LPUja7ZeS/Gix+IIKntbcbNShIP8QO0iRgEv6XNknJng7COUHT7Fgs30xbBWz
Lnx0/8+LuOxiNjepwPuaHI5pEaK97rNIGirTzmKl1/HRKJBtBas5/kN01LInuFzJ
5075Xs6z7Xs/Q0zinurBQCjTzJLKeN+IZLBqzCye20FFAWKVBNbOXgokExTdy0YD
IdQjGctJZIhhbh2e8Cw6L8/LLwl7saXRxZW8js7hZKaF/NMxiMYr09DQr77MejQw
5jo1m9FvNfbmENm8kXb6qToM+leoErSobq58avasIjpM3ywItIOvO7Xza3RpasC6
akIDJ/HGfGc0bP2HsJIVbGCqPlsnoqZjIoEKJke8r1IlrQB6iQQTqf9ABj/Pg3/A
y27mDWwBPhcWsI0PRcm4fUKYUrtX6p3MEIkrW/AVF+qTryWmzzq4zUECTFiCWXiE
e3CV4nUg14+/nKf27ig6Ezq8NYCpORl/cwZ1/N3JbiKBkOvOTBrE0e5+VQ0R8n8f
gVEHerUk2Gj7toii2l0/3agtlx+0P5mEDUUTujRD8X+VUUUxuuHDhQbDyaNANgbd
+CiYOXFsBVq8EHva0/HYvkWJAlFflJHdL2BNmtqMxOKU6AlJeOE5+xbtXl/lN54e
xRI4mYk2AZMnmHYja5qYKIbgR4M+0CHz0cAEVpyP44gj9pvJfEY29oVuceZyJ71Z
gBm8+oqk5ZdD3tGpbCSyG29hsjT0sjaCFyqvmyT56KUu9gaU2ACWo3PwXfVaNHiY
xJuGTw7zwKwcIFss0isOEcaGS7owpRUuhbdqJtZt4aAGQhK7wmOkgTbq28FQJQOO
+QdRR4vWt1boWr0In5Niz9+drmaIhq5PwYi0dJfZwt8H+FF7SfjTSkYyeFsKxzj9
X0jptx+qWecB3bExOOA92mnXy9HOKvyada07i5w6vZRA9IM/TXP5aaSy9hPp/JCC
F+izjDhGp5BBNezytABm8Y3xFi49dG8PWNY5d8m6w4d+4kNPNGA36YbO9bVVko8K
IlepCHzMJRrLhDr92M3ien3YzNaKabupMuIWCujr5iYYO6YbGRgjxR/5aJps8RxK
pLX1nwwGMpQqeEFCZsjkzrupA+mtL4/ZRherCWiA+Gc4wqe2pVyhVKO0N/3IhcSk
apJ1ymaWI3hLlDZaCQoN1iSgNyer4ZeO3PYdZ/G79ErhfHHuSjzKhQeL8MnHnErh
rVv4WUrKQQ7hwV+DuNYb2FgKDw/1EY2pKe00Xv3wcuCcI0eFZ16U9y++eKbzO9J1
vFM0ZKBCGzyDbe1yhHBZeQ/FNN5pOpzLuTc0tz8Ox5pJ3b0pjgMwL6tsMnQmUBEE
SWWmMjKaItAzCIk5T1b/v8p3T5J9XvPCVw53ZxPr6/H/xO7+0uQk4TQo7xpcHi5U
FObYyod1jmMfH1jarCYWiIKSQGbUaNDUs7w44g6ZJAnV81n0i+rnalRyT79wSpz4
2Oh6CtS9vtk421jjmPg5Xj+njWrfsAfkfLhtZi4ISeFUWW6zsKg4ReNPStCwXS08
yJbCa4HhyALI2sXyRS1j+U/DgVfsNqFeErrSAyM1+4Al7TkNDG/ERbpWLgZDaFhQ
wNfV6hS4PS/y/7MhuOfskDb99pHoG+xUBjKRJKsXP6MYKE1iBjrmvwUkA0m0jHHT
KMM6zq/8AOOr7VN16v4hPaqrpLJ6JpC2iI0fize/L8VJiIf37AQhlHds9A9W9M/W
wj9RMf7LZwNx8pkUROP8q9DiI2zC/Jx4P17UZez0XaNR1Dv5WGiYcXzJuTvO/xM1
F/PNw+aNonz2n4tKg3sQLIb5FQLrBM93GYNT7BlSicEzFkGugf7rHcFlRcvkrpdd
tFxRHs85k6C9A2J0PtiNsO3WWBTjJxfL+r/8Phw5+2iTD8WRNUoBlq2RLZaktOeV
b5407s1w/lzTRXAE6PN7aHK7cbg79MTaoM6NW914jUYU4p2u3y8SrzBiXDhA7IUP
Uo0vgDSotPfP3DECSeTKLQ63lWx+h47+QA3WIQ1vnre2fobU/E95/eAqqEFnlGok
b5QP2qUkMHzZwPuB1OFbm4X+CuqipYzWukBFSmsPZG2tJS3ZIunrYsI1c0uPR5q0
9id8p6qGVL9qVhYmwWR5ldwxv62lH38nym+a8ZubCqB7Bukq+gjrDrMdL5TQ1pQm
10NmXTHddeJrS6wWfYOEtKTnXf9sgR5AEk0Q2ZAj4XHcfLJzWCqpIqjcuXnZ+2Qw
9KQ4eOVG7FUxnAijYeA5rpNddUo/e2nNHbdbnxOvh6Ypn2tswjjffE3eMz+qET8t
wrUo1mQkDBxjoTrpK8yyyzFaZd17U3lb9zT/ROqIrh9SaBF2sXR1GyqVf7Oz+3WD
Xy0ft4rAvQTqpf4Zx81vZRWzYKWTwzfYpSIV0p29vylFQujN2gb0KFIQFpfHhPeA
bzv6ERxJhsdPaxHAjeYZM3KiUkEvDewUgE521AFfS08Kzg4CZp3sL159Hr0ow+PJ
Sj4MuMHyZ7W/S/qjdV3QVzIQScEcFKFdgNO/kN96O7U0eXjLKHDEHt+YXarUeVj/
s54eZufLGlkgdNWlfM25YiNYINSGE8r6PmY8TgnJFACEIcVfwe1x3L5B9abwVTVv
yST27V/lcOUT+fbSoyft2PkpQC29Kbh/sgqlm+ksBlSx1R60hSdXWu6gmo9Njdlc
XdJyZbtytyRo0HVHn7yC4Njrc/Y4iT7abDc174LqmtTSydqYNgAVKtEsW0kEWBIW
5khuPKXMgYA09g9JHaQNJWZyWJUf7GOF96NrhV5fKCYF1rB4JR7wUHCGwuZaMFZO
/V+4DlXbRMAR8Sr7tm9Bz/FtXRcV5U72zpHsD2S/uEbs6l+UvsvlxDQDsF4YsdXP
OLWUxvSJZOGI7b9r6Pc13lDQSGqEBRwcgw8ci2bgTgjs0ac3/FAqUIO92CCDrTtU
+4OBbaVDEE4c2EPijBKt7ocop2v4nPaWQQCJiqhZ3xHj0VN2igivYexVrxtTwy7I
RojotJgkF3+DLrBPsnfNl+/kFGc91ZsvsFhoL9RR3nPFOfzy6jP/dCZgfpUt44yP
Bg/j75OuiyMBUfb1EgPxPI4Hnb4OPCJzJIlVWsWNjaP0wvIrTzJP56nLEQxu5I4c
k+7Q7fLeSQWXiynWebvqIvRwUVMUMQl+NcFltTqsKuPb4978s7mK5pojUVqCqMWp
tkKBCd4yQtxDjtP+DiMC4K05cDtK8V1xmp1NhXC3EMRaLAtyEFPsyoTYC/tqmBX6
gS9nBoRbzm1BJ4v4Yk0ycyFn90BVxI4dt/8F0Q6DJXULr0J7PnpJW3YQoErRG/Tw
BaHKSer5qpzuTmR0ZsoWPTCnShEhiHII+AZ8pvAqSqHA+6bDLeF3KtVDX6DV6Ilz
Yhw/uxIiY2hPy74700uepp0mj7TZ5U55t3i6LzOyCIQ94XDpyBBGqfxYU1+Wm/l5
D6u3pzEm6d7+VvVAN4cVl5qIw+9P7BN7n1rlYRDqyLtYoiB3KF2KeONihZvzOplW
vf6dOITxPz/TEGwa5ajznlD1qWGuK4FpgUCjMfCRA4xylJQslgVODv2Ps9n3ejDo
6G/SFVxpF6xunnpLQ7D6A8sQra1PaBtLEE2UL9+m9vqpoquSb7H65HcLgjWvBfFy
EdLJaP0k+2FwO6AvR4uji61b4YHzUO+IU2gZSoZTWMW4RSX43IGVykJHj9ml1IUa
fXhtHziofKBMwWlI+Nt8qPzSeJG/Qlp6kFsVEfw7wITL7AkFLiHfqjT67eYfg/l3
kYa1wzkH7ursBhMtxuDNuWV8gI7NcMHClaxxsLtdUIMejBrmAxP+JgpeqbXtACpZ
4+O2iRVh/8vvcJHsyHu+RdNCegPacPVOjHJOinWYndv/+vXgIUcR94WwM4T82r7y
4BwwwBm9riPapf5LhNfTxDEvZrSo1o+9My4LzeWG6qvgOQ7ROuIamauHA80Q86lr
HZbIZd3Jdq4im9k3EQvKeobu+kCVUk7m+8yAhK9ARqhtN5zVPPbiifhg+1tXYCEZ
ZA+L/88YG/6AKwXJ5Zdp7nE8KlpVACofMUF1hEBzTnV1dKa2Ito+V3KYLVasMUuo
Cd4TjOJT+gvVoTrQIX1YqI1VJEasbVj7Wep5mq3uw/qPEIkTSt0DQiQhx1s8aRx3
u10AyX+ygioRQ6rnZsVk8QJvqyq/giKMx9Jdijbmi3ea3FOEh3OhYR6xDmlJvrhW
Z1aHRU7ma6PiOUdyEmRJivxdXjcgW+wrGHMJH2n2zSx7I42lqYO8WPv0NC3TLJKf
8eccKkoKIH9UwBmd3wzmIcPxkWZF4+qevSqBUoq+6EO17yRtVfzaAkfDuPQJwxTQ
nwSQFl4Nyr3A6X5jNgJ9/BQnKKvoB/OqmUEIvB7Dd2aU6mK5QRKzrrMrMuLWv0Xh
hnGrsKmkNaQ1kLwBSdDIrCnLB0GDgE3n4DDMhzITyCi/sdUw+C3CiDeW8GcUFHjN
ZiEP73Q1nveuuhWhBGZd2ARuRQEFXurHP6qgbdJOOHrTwQHy9DDccFuHTN/fXo0v
cCIAg3EFFpZ8eBoQtoao6MHQZtZc9NHk8q+XgdWESY//XtlxMxeThdV1EhGN/3dP
HMNwyJ9OCcPMCWJCz2+DM6a+NjN/G0IluSkNfo1HUd8NrOCbY0KMsNxcN7f1zGPX
IB5dNSGenm3cPZcJqQ/45nPdRbRXQ2hYICA5YEDoYWI3Kssats0CUmicqc0mlSqy
DzaI0q5Bqc+l2LnMWC0f7nazQGHQlH1sS9c/BmljQhsagLmlzjYxSASQdZobX6WH
H6A2x0NHtreSvLsDaoJuZj91gfXYYWFv07KNeb0pwcOhMjXmVDltqvTolnwPp64h
HLI0PX7vYa6CHxkdfbv+i6qzcB1z3s+NJJPwG+ENz4xfdxrbSTcEtO5e8pjVqU82
WE+XVpAyEn+OgdA6+IObetCyy+shOKAGt7+kNHhTu6YO5ggA6lb3Pl06A8iCR2/U
Ahsy5kYgJsys0+c+OsM47MJVZYswrK9c3ltVpuLSTyAF+G8E34Rl433yAfFEJ92V
yO9EiYCQVyenDFCgrzpc8xQ69IJM85waOSWkhaTrT1k7EOYqxp01cuDmuG8nTSZv
9LKFibh5yxXKDadPV07QKRgbDHedsOMvcQW0S7szkBXFTb7+1l/z33+qp77oZqk0
Z0rCK83AU4G0uY4sAVj/cYcqRkXoH2cf7KqI0Oyjc4fSWYR5Ytei2hIACSsewgkt
BJU/UeHsp1woni0EthOO7928/gwBm88QJ/ihbFnxQnwgn55yic3T6bHS5GUgE/iU
WTSZmffvroV+6xoFvCHRHnmX7Z5N9tC71gNudkOJWqFszInD6OhnP7SDO3U4sbDk
uaWhccIv27iqJDTTU/w6vLrCDTnOewdBJtjq+aMjhKAfc87dY2h/1yeYNAGRijS2
nNEAxd7CCmIuITMSkXobSq7y63Y2BQf65KssgAG2gsSiUX/QU5eNtbAXZ/p4kUEx
9kElX6wrwohOgZ28oQjooRp/RO68SOy6Rlzbj2w/LtPpiREFrpPNa4UeeZy4bRQ9
BE/+vQRzL46icBO0SO/eC6OSPtYjaVfa+oErxmJzPaP4NAwUOaGAqcBwj8NOsTG0
sqmthMRbs77sqxmjkFw8dkiffGTYXVWlUddkxbJ98//ZnGlZr2UJJqmNxg4Qd5Rj
CurAhHGNwsziqKorB83+O/lHh+/nuUxnxfGSBcZ3chmNBrFxSL5Yc0HvlnRNMnRA
ISuIUggr30UrJWege72AkG2O6hOgmsaMR6taRN03uSrQY3pmlkv3Sf1p4wW6N+1n
Ol2PqvtfhVz/j6gf15gNsmf0y0qf3WkOFXDrtGGXeLDz3BhpAOTEbF4YMocanVvA
svaG9FfRhxU1fNw0DPhUgj3lQb6D/B/LxKAcnw9BYy1OuiusHDJWTmqkyfrIgbyS
nTsXTqb+IoJXx4TakgmivJY2HXj1ZWfLbNPJsfDcWWKuztJleV5LXKChQZK8/nsJ
moPIl7bR92JQZJj36flIxLQD0NYTOOceUlMrZIhXtT7MIR14Q8c3uyLMCkK8JIbb
PqkTNtLXg1l16jUgh7PBCsPs4gupSd5xsuxQBsYX6hFNjheXvr6iHRvc5cxom2sY
eSFmHSsk7OZ4SgJof4LfrHocWNW3+vL9sBw+rkt/JbAlVrwoFl60mP3xr3BeygIm
cQ2ZSIFfBlFgfQK9swoHlvoNHNL9JeN+js+SuhKcYDVgPUMdHjLnISilUQntWYrZ
jj+Eo8gFG2XkKvM9ZhhsY057IIVJ9zL/B+qp82MZrQPgHmNhKhB9U+43M3NMXqcM
l1zcX0/V9XGQxNq4mmDbR2toIst6bvsC7Ft7mbXFdsQzsBFc4KVA5SsFFpDNSD70
6iWjv74UHllic2cO8Qt01iG3dhVP21U0knRFLnVGNXlEYYGKxpCLo3rVlMjuMLk7
RBq7yNUz8y02eYxuLkrLqbwxc+RZi+I86SDCYNRDHf91gT6NgMZdyfCvE1fKVpc3
5KtTmH7WAFVfpPHY63UI2QkkjznkNyRZiRNDaH+3p8KteWcLzkZhG/7CfhdFWhyC
398K+xqnk/pSaySB9F7uGNgyyx/wRnUlfztHo5rX3Sd1JxGcZQOnQiTj4tu8p2MG
NIhaBkKvV7FLW4t05TUCSFOEZcuLZgKujlZjBJ1n27iI/54lMykm0w9mINZ11MmH
DVzfQO3MA1kgKPJVr/bHge8qU36hLs9UY+tS5W/Hol7dHAdUQ/H2kmNy/0Z1YfYv
mmlzmVzSQ5iaBDwq8G6Y6bLzHtZ7YL0j/pBpr6UdyHrZFuyW2nCLVio7birV3nDA
dQExf40TyewvUtbEigaqrqcSjMGnBcgR3E05i6N3qeAFIhPu+0QQPe3fbjxix2B+
42fdRNhcy7PnNxk/JjAM9rQUh2JF9TwVBP8Vi/jek6GumrZkhHMKZ5nz2PxSsrKy
eh2/65BDQogbyhS1xNZOqu+VlHF4RKQ9W8Dtmyl3YpNXxCuWxe538Do2VIcUUHwZ
Au5DiiOpQNtWZinJDBG1669Sa/dt3Ygtu2J4RN0ooAOVKK4Vp8cITSkdmroOxwqz
Kh18MgapmNe2isGR6LPuTcBzkKbfT5yixhFtgkoGzr86gqCenojUNquqhaHiqQTx
21J9AhKOEk5Zm4oTQPW/BmSizPiMXggpKNFtANYdToyFtPUDUtx1Cgqkq/mg6DoH
pOWKlauxb0v+5QftvC/7Dpo1BHlJveWNS/aTpD3mE7Eq+Xt5gwAtcEfe+s0Wbwvl
VaH2DlzSLhIXNcYgxrcZiIrN8Zz/T/27zY+glgQZ5balnYJTfciZI3L4C9fdRkfw
WLAurhartKrnEpHgRxrp4YRdfqr4GIln6H9hbK1aNqEn8fPd97SvfKLQYIhMrpiN
2x9IWsdIFIvJCE/s2vCSyr1OSQ1fgSlxbbUKbtaGFcsS0Zv4xXysV7NdD/wgj3up
xBcAcXslZzyHMZnzMXEHKBjxvj9MDb76aHqx+rxci8hmz0YkIytAhzXQFuyO5K2+
0Gd+YYBm37OsC0XEwh/L9wZ1OEcA0Mi887OM9jfpE4Fm//XewaPrxpG1090EMn2G
v67QJy2K7eHrqmwTI+GOymRjCI5zCnfOrLM37N98CvF2ZE2+l6ZnSMnTqDc+oj/4
i+11707NCH245WsTFCyXHV7N9l7aIW+xN2gdT07W88HjArNiRDyQKQCNrIptxTh7
hzn/wYUW6Hcaabomu/c5qSof9u6wMXVTMniKy6CUsHEip6yYwy6FpMKsBjVzU6qK
FeaYUNJ6wJ8fL4aFDFp3pHr8z71SrGRbrPdUhFaRI38udLIi6iQB/xEbn0cl7U18
s4iecgFaHGgWjFD0Y9s6ynHninhTS09ATkPdy1dyr7sm4nMpnxLRWofYVE74QOjC
5Yy/lplcclu1t6SrhMg7aXvwPIIDtfnjwa+/Mi9bl23qf07CMXrVbCXVc/s1YXfj
ZOyx8vhYz1JrvgWzDy43p2LLgDjKLjjK6pY1a4MSsErDDHtYQGXDU4PDkDGwX6Vt
VENh75cm6W+gRuW4iShMrgycTszPnQ4bM0VkL4OQeh/J7kA4vRl6NCTkSdw64BXz
lPZ9BJJ9wQgf2wC6TgLkJILzagZQGFY3df4GkpReU1grtru2DdJV6jXHRNn5PwEn
RtMER2DnW2GsjLD65TZCm08D4e5tSyLv7qPUVudhCuESMmTMu4DCKrcjyz6zoMH3
K5RbEMcBvRCta2/7UcXf6DxS5OIsGDCfkg5OPd7xIvz5mwoM7hFJnUE2+T4H/2OH
+btQRE+DcWwhP6g2AfboZhRTs0p5qGRutkF+T4ESUWxN6loFO3tMFJsovgUtKa+V
ji0UaaHiNWUMvmClBpQ+XIAQJdiE/FboCuSmthJrQ58UyZlGNZwcwbxRqdhLnlwF
SATnsUVL+hIT6DejawPNF4w+UdAhZEzfwKvZRP19Y+zFJfte4ZJke8wK6RYplDIz
8EsCBbIXxxXSqylCERdYk21RMdNx45opWZmqzUS4r058a01QPNrd5PZSxmeEu1/a
iR1yFHVJ9ZIStnJT6bJjYCDgdAsyZsTVuavmYIW2J80LeSOsM7c/EbNdpcLEWZrl
LQc29qDEuChxbyrr08Mv7PwONQlFSC/NohzOEYkyyByiwlLtUbO53Ivz9eIs61NQ
lt7xQorb5NQxHIKEuLo76WX//iBSv9VGdravD0OTzkIO4Dz3bCU6oDlMxNEVbYvU
2ywOtyA4uTx88ZhtsX+Yz5q1knG2sFl/Vj0pWq8KhGlf+uNkM9k/OLHfNcoX9tJP
yYcRIDFKwIstr6X7XihmxLj9jYvjTN2KeOelVu+zKohpy6KsbBOLYaDxd0j795VY
qpNsyjOWvPexbpSaQ/WT/3NyOSfMT6U8z5LVJj5s3nH9lhmJfXbyOzxcTo+PX26u
yXnEKf26DAt1RHzuk8/BNqZdtl9UmlhDOaxKcewUqW/A2ctdnn5EKd0WOMaeCKFe
pEXyQDKp8q5HnNZBSYfBVAmfT/+5OQ0TfQL4E34VDlpZLZfkRoy9K1ndKLsWWnim
tltouMyX8UUeVBMjmWWNdZ17ExieNdhsp5Z5N2EMTl4W5zmpkULTeB3pStTNooBn
hwyRmjI6tU17UxM++/J8sdMjp4SaSCfSooFQ3OkM+AD1ID2Rv3B+JgdqSxjRQQ6v
5G+IL1vZnebjbh3llRbFw/xhEIko9L2H6wlQsgq0VrmC2fCUiD/OT5ye5sfEGLC0
ctjb1cUsq7+DI/TmigdsVn+y/brxzqneHavCTIru7SbA57h7UhcuOazXPg4xVORU
QJR9vcpHOZC8sU4UD9jd+Ice80+vymYFojNd4pe82An6/kzSpLeCSwC5uxYvZr0m
cb2EGcY/5U+Vh+XFdhz1XzBCozkq4TVZEV5XXIjj0PtqxHblDy43ZM5BLm4/Bvs3
Ju/d7WjJ2OUMfJ8/3JeXB+AJ9t3PRiAv1RLkwpjhVEfz5e6rpyuIpLJzFy4sfprk
Qno2Yx1XgJ0HsuGbnyKc+qaoq9/Imm4bOq0bAPi0PPMB3iI2yzA18AqWv9hs/tor
01N9SeIsdYGgRKuH15zrmFZBNzp5VSfeGqNRuHCsEPxIkVePJb7k3N/rFpiwG1TY
sDuLZYoiXxle92hnbQU86f2xFd57A5CsT3jwh/epT0BX3SqVO33bVRuiUANZN1GE
ybfm1JZruAdU+ASXwYJ9T21TCN6M6AytaW7Rg+YxqBwsL01umDcm/xjXgYS0BPt8
OahiuRgUju2LRyBk0gOxIyimQAoIDrdiYbms8d5peRX57HlwbhEEL+TSG8qzvnkm
lsFvSnOLKHbFXJd9p5PDA5X7jom3w8FBUFqrx4Leh8e8jRqssYKTgc1AFiHYpg+1
+JOEbk37dbJbnS5Z6oIMwR4PHiiBFKMXS2rQGATMZ6Inl6Z3NRyR4cR61MYK/Jnh
7A2KePJTDLdB2V+jNQH2sVN/S+PUnwHTVqLf9fXcvFXIySN+E5/MwgxLKnJj0T6q
W2B68rL+A22WGERWT7JIYcOd3iQyEIt7pcMDrt965ry3zMwnng1dTCpr7LItaxMP
+FiIwNYJBaItenH9YZH9FeD5aVB1NFTqUz3hB6/STHhiK/yFcChNXg0QpR+v6C2s
bnenZt2TVhJpHATQ0D/XtKB4S11F4mvTc8isStoeKWQL2OMYQkkWxjD5sg7AHcaz
LADUqwLttJgMNmV8yJctTCoaldCJvBPUXSJBFJwUbTUl+mOQjCW1QYnjDYgHKOfK
oTRVH8CicGIBuPcCOz5r00+jT0SgzQQ7f8Mkbqm4DdKOxrbtbphmt8K6b/5jf4Za
WTYZwGBoJlFZGBOh7Yf2O3VEY34TRXGfamEoQHLvivhithz2ZAgx7JJpMqzN8Cjk
JAJnQV1u/MCMlyrcBzeNtIumQu8NUNUGI93+bsZKsipEpZ3HZirJnf1/G9W09cyQ
GzuXTPORixV+TyQ62mGSwZ85oO6f0CtHdSs4CRWCKB3Rs5lQ3QX7cmIj8zlTMbwC
OUcJB8Uboe/2kHUhIy1ltruuTJiPwjYG6fc/N4xpDK57Mn6hWNwpo7RrFpBlkR+b
6pYqdZPgTuZ12HIRgHrWVSOqRoUWTFfs9/TFUeTYFEq7znNS6u6hvJ/W70sglf8l
SMkzvcTd6/PnIWRtiOCi4WkzCZb0W+5oLmyea1q+9fCJfEd1tQ6KEG7WvzKjZyxP
6Jfi6VyXFJjmfEY7srTf1NZLIDnax3stqXel0jmJDMXV0dfDtf9bDo7a3zYwv4RT
kCiL2ABNYZg1XfQg4TXI69+RS/9ygyed6xeTCemwZeJidDVu03dqfayznHjyGZWd
MuFk+i9BeDhtrm0mGea+93lT2nRLrvUeXj/uN8P+CvcaPQcSYFjA3ZPK9ewgvowy
4qwokb/VrEeZCvKbeLltZPbDUl3emkQLgCy+cInO2jWsW6nq824/JjC+xQ7YZXvC
WRqOKKovNNFjkxE/WERssc5/vJkqsGrnC0LEzxReHJsn9ESLqEUt5QypRIC2OWRX
cHVSMELlHzbrYFg75mNNbLn15ttUaICmfxJO89UsflLU36qDa5HVbYEFK7a7Ntwb
HeN6u43c9jZ6/fUg2x5N77LL7eTNCVj762GkbE6pXsmvSvVP5be9znMQyj6MRf55
tfPZRG+GmIaJhHUcmxetPRlyZQlzhBkf2x/KecFO6UjUGkPgDeJKwRqgnl1lwjdZ
zt74rS14Tug7/vOkuugFe1epeiN7cAVh/eppRUpEGivCDjmFQIc0xcoKInhhKARM
HBLR12g6qA3AQ3VO5Lka0XBQsaCPAmuB6Fc1UO5XSXf4XqtlrGLUHeUCpmMHOq5h
1qRUIpr2qUPqdWoCDebA3WYDpdxEDpsqB+eAnAeCUmmi/3g++mCj/E8ZR9x5lwjo
xMqnFUqdPHuk5DQYcblmsa0ncbP6jRpD1cQ9bqTk8BMSoFHkP/hwK9AEXiDiokgn
9hGYHBwEDKYK2EvtJZ0jJG47nOWP6m8QKhor7gNMUsQpaPCV8e6LEeAgjm7CRfMr
+q17SN5ESkJX8bmyyeZK6al2N5EUWLtevXsNccrrInF3u6eA+flI6qiFBWZqx+31
aoPAH5oJJnpag/hCGla2cZwKEz5UPvu5iBhdMhIM7sAbjAFh+h6gY5oejoJclJQf
22gSvrqW48LeDJ4PZgI1MTdmI/E8Mw+d5SaKAnGcgNX70mUiuVvHSWF3L8E+wJjo
c3J4rF5xuyGytFiX8bRDpnIInFAdKj+b2/MuQUCB69ODCE4KbeFKFq2VTK1Zz8kB
Wlf+g4zmyiN4Wm2iO/gb6EKYraDKaaCg4a1gZXYjC/xGvPugLihvEBjO371seyRE
M56NCcU3GycxXoQudF7Ndq1BkjGfucQQ7E736hmdb5lp/QElqGtli40UX3/yo3Pt
xEQet7laejMf1FETznTYNcMJoztAPjySrm9yHGRZ/7oGeSlmpuJgnrven+w5xqAq
eYv7cqIeoe15hs94gDDyWjmcFArLyZsAEtNNBoAakqZVt6SISA1b6rpGXJzZqfBu
N/oQgVRzelGsG3g36fhB2/l2hmwLXGtYiUMRJedL+CdSqZRaZxLh3+an1QWLYmU5
hyUqiJBNCMReifVSRurerAStI58Df6cPOZa3G5SudeMMJQ4jvGz1kZfm8Ee6+CIP
HJBbN7UBztD+to+5+TQLE19SugUlATESlPHqyXpTDPVQVQXcBgQ9i+vm8fjfuVFz
Nd5hXxD7VeUAAAY5jsp117R4rGLU6GVbz/kqzAVCVTlT8sD42JKKXwFvy2DD8bBZ
dcqe/dIcj+FDxth1lvjPhpLHyaGaAO+AEtJrEGrVN9My5w9RhR3MiLYI3EP5UWC8
AjXnFq8A8ATVvhXvB5yT3niflmM2Ovs73juDtvRBVsEWoP11s4K2WiRCETKYPzoP
av/3JUYpLoptCTcRAID2sql4VZsWb2NuFV4Xt2hmLvpmgHecbI6/DXkzA2IGjOoh
mb4l2LHdHku1dQ4Uy3jtxkd1lgu1tV8ZHgpyPcq2Unzgv4fnrnF5loUoDA8Ag2AG
LKwUYUnVx8FKgihTDBFrD278ftdiG2emJiezhzhsGFUEEyLUga6ar9QbPPJsQDKQ
C/l6OGJEEz+PNkr0bxFXV2C8POW4Z6VYPPgmil5D5lVoX/hsnTIHhai6MlByo7ud
Rq04O5sKkPTtbs9CxIEsxjQUhvZZIzGJHDXFk6sN0iTdVsG2JSxmjrpPSzw/tYyl
SUrE5iRQQALXVmhdOAhtvu3VObAOrFkX+RROH2x+LJMg8fDwDxDHz+R3K9EiAvHP
Gim7caVtiCsT+hb4J+BaQ9YtOQsAKBhr3xfpUG92Jn0nszU6Oi1qprD2G8WsNlYX
FdA9hauv7btVeXf5JzOXgyytI7SysflyRLqPp/7+WhiFX1mxDu9+oQITwokQMBnv
vVFYk/Sa2DftqM7xyD3XBlN7MNBeTXB8exQ80rEjBgdURzu3VfeLCWTmwVtuiyVZ
LX+5qMe2M/Zss1AEpShudlZeN1W+fauKCcdH20DQX5ll3c8FG9Lnlv6dt5LQeZld
HBm/5lXq3vzsfnbTsc+tMumDUXAsP2bCfYRnBLldx/qF4irDTulJYooqMxi63Pem
Scu8v/AypI+LjlJHwouABw5Qd4Gad7V1OIQag5Wl1dFGzCEGLzAH63MaC5Qmanrk
ZONzvjo5jvquORit7DF4P8LFHgdZAig2oqoJCBAILMaAn0p5B6y3OINiY3g9TXST
x+1LH5ldjb9SGapG6gAdVX6E01mHWGdOhC0ITz6NN7UeIEXzBWgVuXiwWUfJ/1bZ
OqAbO9xxwuC0y7E9LgYjOqAmacImhgDdCJc8YXAlWhC9Yo1ih53hI0wY3XXL7JDe
ZDh4B+LP9nMyqv/QsxC0z3mLFFKO9ym07+uFGyOqmzc9hfMMzmWeI5cl+8PUdfRh
pDCg58XIxRwkJMnt5lnLkEJnWL4tyRde661aaKWL/gqpi64/RnEOxZm42NOCXZ6e
ASsNnrB3c447WPOGuaGGvzbqYXaHk4C2i1HsMNXv0ahRmMq+97HUZ+JjPLrFbsWp
S9675v7mPMx3o/DZNWtpZKR3yX577owXfRlydIjbDwYyO/YETxeUu9w7DMrZyOgM
h0yMCtVXafLPcT1fVJi0KbTceB2uuF51L+47FveI4zPGSYdjE+lLdL6WA3xKY0Vs
re/Tc8nmch4xM5I3LbaRiKZbHT+qMqhWQ/v4V+S8uQTtX7s3ceDT0WNvZW9o97EI
4hCuDizvdXA1cIzFW3lpjLEVYoyQpZDQeHR8tQavEv0nOZtuyGAa9fEEkqvmD0lH
ent1xjvIkDSPZ2qp3SV6gkSwBKn5F8GssCLzKVBdqiVjwgqBoQLz1Pn1+tMYfpL1
JjYWRCcq+FGv74B7cq+T/2TVuIwUCGcEsJiOZBuTEuyHF2T5fr89AJLTDQNZatzH
Uva+g7Szbw2RTy9SDZaSO1CYBDBFPAkS5w8AMZ4Lo392dbTBu1IBBw0frDyPRUiV
0ocJQYyW3SJ7wTwqyGdX00RN4y51z5SN9wAvWjsTIbjY3PDHb54mjBgFkWPy0B84
EQIUkHW93XTkjVJAHsC8ATxk1Wbdt3rcK9orGzy2OnGf8qTj3b3ywgqWoeSRQn07
Pu1sBD6/jgubd6qvRrBZNgmZwY2Qz9+1JwXfWGZKjbuV2zE+2b9O7Za17P60ijYg
ws9CXS3YSSRFJQyNnF3YpnGL8FvHvg07l67oIqv7V2IDlEB0vdlEtKIeDSH1kaTe
8kFnqbg3C3KaAZPuTkJfVBqR1YRV1dylK8BmHnTNqvOxXsCp4Uj8kMeDTA4AahIW
+rla4fnwP+VcJjaY8pzebYHQ7Z1eWXWuTPxIsFk0+aWSCkJoB6W1pOpoqhoPAt45
JTioe0ra8q74tAUFu9FgnEq4bbiGmuyMjA6Mte9s6cIpMy9P1acnuasXM/rWwKMG
GfjAgKYXPC6Z2LsrkNl6FOcQSQIk2gFPtPDLHXcZ8k+iSSAXqn0WuQxREN1IBSG8
NEan1zFvNS7gpHYCDU6hUDbzzcdtMSF2nNiCe5JuBSMkgYXmH9VQStVrnojJ0zHH
HTuMA7DKqpS4ehP71n0aXoBpTF0CKr12vcshQqIdKbuIVHNFNT5cHkAD1QQmQYnU
IN/Kndb9xEcZaLDxVJlGu+I+bMKbCQUplitbFkEuLF2LfXtR8h2NLIfebarSwIYT
gZRw62eeqCIqfqd9TDax3pHN8hkJScTIr/9RsoQoaH6hWfv85nTCkyemj4nHe9/D
i7ROvI2E6EQJ6e5uQdJz4bvXZ/3M0+bD2OWZysn17TZg38XaFHc6uiOD2QTXflDT
C8yy4jxgrfvmgYcplu448IloR3a2/rLRW+Bui488OXC5FzcmBR12iVW5vXxQmbfA
HMBaLyobLsO1K6fm/ey5HwERwwb2EnW10lpjGYYH0GD43iMriq4SQMn4w6Xi+DQb
AYtBVS3NXn55sBrIR0HLxEH/ODAHZtuRisbHx9zcHyHLOVNMg1OJG9TxZxRneHZa
AC0IUNJfbKgZYA0/X2jz+9Xr/2UWhzZXToq0g9VfhquRBEXER8UsvBO9GFHCSKp0
1+Sh76ljjbLszMZVZtkc/VwLhRV7c0DdzEOcR92QODbkdHX82X91/FAUoxI6gHsN
YjRspRyNrdz/nYy+V6mBDv7jUd6YkimSgPDaoPxpDZugxjIMvzMjfV2x2LpfB62O
7TBUZidOTxzNLMAN/ZpzQ8vHqMhtQn3bleT3uG9FLOS/BU4T73KD35zMSgwhitoj
W45ZQT1tdk+N4usiB2k59TMGvwE2i2fMjC6MtVA3gWqUr3DVXZe3Nb8w1ze6LpFm
7XU1ugjgznatCsjvdc0kZC4rb5b3HNQHN7Gl7pOpiFFyvCiQfoJHxZqWqie5U5ef
EwZ5Qjl3jEXFvHy1islyS9N1ssIMvX2wUrctGfpulWITaee31osShBq2EFDgMsct
Wc6dnHpUec0y0lNJ1Dr21Sq+BTqQcGk4UPY09L3Fd+eW28dSni23YKIKF9iY833D
w4bxBp0NzoUJrtHtmETOcmuldJDTXUaeINCR7kGGhP9jTmLljXMMqoKRFoqscE43
iX8Om7EDmscSEEYlmC73X07odRFfxx954d6+YhVVC3sk1dk19xHTpFaUXLo8vkGA
jfDyjUX9LhWdXs32ksMrXApTY6cAJtplVikEdCUM/ObJWqYlD4h6ugDdsvwuZhBE
KKB103mCu013nl2CP4yt9VjqrjYgTzkJyJXTneA/V1jINRDLMlWKCqZ2MwOUqWXN
yBRVtg5ooirJwzqVkwGmX805kO59uyrr5o8/SMK56k4O4Jl49xnYH23dTscOotOx
fdqxPJ4kKLJT15k+TnIFgBwqjVdfn0sVYvT8KYuwZ6uNEq4sx1pOy58T0x3Pb4CF
cDE9ZaSQMREVdamZjYcfsfJct98iKCzOZnYSw6MHTuXmrNn7EL8+bOSJP/c5JVxU
ZAxFSt2g5gN/xAYVpF/Tniom2ZhYDOz8doG8TkuaJo2vNatcWLVGw15PoYz3oXeA
VbFe4mrA7dxa+Z0qX5PTBXH3K49DG9sYY/BDLSE9anw4R8i3m07P3Swkhnm6aYRr
OSrYy+tKREgcKkNt/u/qJ9GwbCgdHZaZw+5IEWQMReP/d+62GORQ07ttCVAMtTKs
mBoYO9LiiGhJgYWI1n9j8N354b72xBWgF6S2SqWv6o8rGqjuxpAvqTovbVE1fJHZ
j8ivzhjIP623zyVAF8yJTNI1hpj961JtaQ+OlrwUbRgXm6vYzOxT7Q/P5wGdR9nQ
4Tg0530EOMWLQT2t3HzW3uh5QXa3dtIa1nYXQrmGD2JdntNMfbLYuJj6uIQGtDd/
ormT/y4uhCt6HTIDJrKAUsuSx12v6Og3eTJnBXphvipN0Y14a+DWf5hR2jFFLWIg
RJMkUQBvgT/FpgjxzoxBIDr1EV9Bgh2qcp4jKWdXNj8klwDw+jg2gKyTtiD1xaXt
GgkYcn2HjuwMTZwnsYxTCyV3P25eceaHWdnpBH2JLOB7gpfho+6SZxsikXWnp8gc
ar7WidoJ2UUhjhZP6S8zjzEtEgJLlnX6LLkleYyBaEE8se8S3tZm1tadFaJ2ZykC
D4nehg3Liyx/O7WlA4m5jLLpzvmnAaULaypAuiEE7NZfj5Ay9PRBGafgQqvZK8Hi
ODnr2UpNU8keMsB46ZUOdalCV1/si6BBbdITfxpCwhoMuTeaN2YMRL7fnEoGl0OA
xcdQ2PvhPzhUY5OYVrNk7gGeOLN6iCqX3Vgn4l/7aPocs+HGHoxe4WpEVAD9CZCi
hBTr97GnEiEvx6XWYOH45nmLRWDj6RBcWYBJzyyZShB4H+g1iEfhfWOqOMloRb9Q
Rd2yYEMaHrF3DGATfCriWRAVkHGlGLAIllBxj3i4rZiKiqnhqX6vG2aPOuA4oEpl
+f64/uMvCZyC11CT2agLJ2dE8EVNORJ+kUDVl1ClN3COzwfydglCqTZ7Dhooye8q
V4PjHR8k7KVhENtZtsb77sptz8nZoRNo4my1jGsgtOjMZTVAhXpzibD6D3jlYw1Q
SNuFQKHk11yZOukO4ThH7A2m2NYGPI2FQcJNjRJsyiOUh657eSa041pLyPCM0B88
hoiJYYfGDbKqRBjcBPCDSUlL8f6lgwNK3EFpnJ4jNR6EX1TXSxF9Qbw0ety7siP0
9QMMJ6iTO7rXTu5LK8E50AzV83n5cSlerGOj+oMw3R9oZPBtkPgWlt5MsrsMezzq
eRVQzz0NOSfMNhFZu9PVG4rTw2KE/quc4mQc8Mv8fcmeqEQXpZW5ybnRy6oZnXjZ
1Mn4m33xBMy/vtOdpQH+xkaJ4osQy1OkmNfktm5bzU/I0OI62iSQv2WjNRh9ykeE
7W4hDruJA/hvX4S83lBKiTuYGgadrZH4UkmNaisVHavwp0g6wnKCGC8IlunclqJs
rrpUocDDIDWSM2g83/p6YyB5JwJ5Vu8pBaON5SYcBdxmhmxum+FaeLCUZUjrfxb+
39R9kxHM6GoVwPeyoyIE7cg9tePPP4gnNPhkanJ4ZMKLMAeqXWBqXNhdBqXu3rHW
MXQO9O9Flw7mIpBVN+IfooMU4BKxQ+59Y6lF+Ja3y6Lz40mflx9qsxBZHrQHGPKN
3HQLGrTbsDKj1qaZ+ZF4BmABBLQ7b5k5qPKureheCMV2ypA/Zmgo/GhPjiby50yv
KtBSkxb+jpMA55HC2Fbz8w1B3R3t20suQX3Ls4KwESkTy+L7h9FeQVkausNYk3Hb
+rFsgjPrjavYiXXSdWgjPG0/RUbkDjcW0XbQ0NqVb4AhDfh5wJjRAxeEGzspUxRS
9MIXwW0olwLw2jQ2LDdF5bW7bxBgBGKOBCrRF6aGm72wuLfjs0YnAhok7eLfW9HP
OfJZhbzqmzUbQ1je38t8pgqdn6C3ZKznNsG/uz2QfMaJrO26KW7Tgvydwe5XKhG8
m519i2qUYZXN3fPdIfNh1AZbO7ySssaB3FLeJuIjIqtXmQEdMdSqe03UpETmXhrV
zwqmtpDILe2ro8ePduRC6uA/YNjc8sejRw0DggQy3veXA+85LumiFSLn4O25nc4L
dSwok6eyMFsRSKVRFOMjLSwNr9EZ4chzkJ+xQcQuGP+KS0/pmFTMx4qL4XmAcBMh
89sMbL+xmdBhlyRXTv+gGCwhtUUbfmeGRrdPwnakuZNQJxxr38p+e2V/olazzdmv
BN+PXdcMMP/C92pKvmJSQNN+tYhlMw1imTE41Oq6Jtuq3WTfx13vJZ2gUiZvwBwE
xC20gd9iaZ9nFPx6K7+AqLeJGwkcf2J0LtF2Mk47m6cLOcMor1WIgFznSEAXa44+
EA2UfBNHKNkQH5bVnNya2W8cF5FkDLSaUVkgzpixVIZivoeJpYKNO366mW0t5VRe
ZFB/AT2KCZS21hKHuzoPYUp5Sc3wB+TQO91C94NpdGTHoADhWA3l2f1stK/4MrVn
x6LXRMm0nn3t5fhFey6i4JLcFYyYP6thDKph5R3qUGJ7IFh3+hgpu2MrcDVYCpQ0
z2PeUCXFnz6Za+GyGOixMFBecsbfxsGMbqytYdCB82xROqGslvhahS7b1qObqvDq
/UOG4hjTD+46cftKQRzrY2FjGz0RqWz46Yil6RP5Pc14aKEALhfcTU3zvVmLW7cH
Y0Llw65ZqrTy3OjzpWE8dbLnPYeVzA8Kq5wJC+5FNwZ8fDmRcjXa+a8FFlstvTCG
Sz7IuAKNBVxnX2NnB+YdVn+M79EDM9AOb5nPbuF7f1UxNXclzKrFrnXeK/rmyTQk
nwc53yRmLTLNMHX8EraFFFXtZq948u7abcF2lfNepbuw1H1ps88gvENqTeX8QT1v
h9HrfFxA93y/sb6XfRf+3ZWM3XB3E6TF6u5HD1T4fdSSjsXtPrN9GZWukysfJ/67
DXtPv0YVEWe3C7JQh3Hog+coHkxjfMcPEtsL0qg850uj+40MDPG7V71pbV4n3dgl
ICe44R8C98Mhig31JR9v9xd7M4vfQII4KJl0tf3x1PVANKRATq+SnIB2j3k2X6Tz
P6NFjxrhfVXNGaFOg6zlbdTViz8TtXrejPyqgb45+uAKliHOxPhIo4aErhxAO++V
JxvD1TkWywHINYBPrH02dXLXV/1UHrZBqVSOxdcBnNgfQms1yTdzDKRHStv4Am8k
4AGldExxLhY2fUq69L7J7b2d405e0zOyvpy2lU9a1xNfezeE0TO3I3UKA3eFdOf8
bUeGCQ1vzLrIyzYR83AKq4VtBOnnMLNmscHtt4Bctr9FazuKGSTcraykLO0AjgKk
TRkloRb0jIpgXxZMTooFiZUu+wmwAm17yE9IOAMw8LdoIl8Np1ujHs29tUVJawnZ
FzQfInfIL7AwNmdWwI3jYJEl7ko2CUZI4qrGRUVS1kHHtPaCaqHjQt7f4Y4ALW4d
5np1DWxursdvgJKRSLZbaldLNE/SMN+dexA4eV0L719vcF4IqE7gT70KgQuPbsxf
k2gLrn/0UaTgjUnNqYOcI7hvI7wLL8wJh4R50A8PwExGeO0JYv+2k1pUbnISx0k4
0/rlE++gkZzVu2/i14VwQZahmhabWeGj/alSgMX4xOTtGXifDb4lKxh05xKou79Y
KvJIVtYXcWG/ob9YDrwJaX7ESFt6IQaM3Wk0QjC8cJH/lhD6/SlExYq+xIldtS++
RhuB3Rx/9dyZG8ObJD+Lneci/1IaFv6k8vT10T5vzASx3bSnX3rUBp3Jb+NFJcCf
J9CdfUk6DqXxpklfe9xWODMZC702mVbY/OnYfAddyVJwCn+ccYPtIniem3qxyNLJ
aEOZI5TVJKflMOxE+XQwYc7wxkPnYqLnhk5tOioB1/GmEbWkmfIWHhCis7IOU6KX
mzD69Kepg+kW1MVZNGpfxpQ3amb+bzY6wcEwu/Wk4i+StegR2cdPAwFK5GVvsNjt
aRI6NeakSQkxgdVNwMkOAJFYzhDqJSqbJVzeqY6V0xa+N+YYUzC1avK5B2T5aUFC
OVGwpaeHD593qJQoqcZAaWrK5hg+YgtdJXYxcqBqJH3s58hJ/y5EFOUzr/NPg64e
GnG1ugDQNQQ7EJ8DDEEjgf4PtT0riVf0nnVkGvobij9v2zOnHcLSbl7wFE0zpS2u
HCacuXzHM5igo6S0GJkBBa6SsEtoCOBBdWlpuj0jjMUKxXz+oiCMEhcWTZ9t4mig
6UAjcz3KHN2al6yyDVNJcE6ZiEIL7Zndn7NL2ViFODXystsVDnckqpE3yqX2aoqF
BzsfBN+e2b9lOce/8MS43lYjlp5uOM48p9s/i0QCPfNQx+5tpylSa4xz8rQDyzO/
F4Za7I7OBHGE0VIcGV1ttz1oxuQH7puGfu8mG89mZ/h/M06AYF32vZrWz4Bwp+Ml
fgcKXrNmJzpSWWA6fgK57IoRLLVRx9c4VJYKjyj98Z+i0lRzG6Z6fV8p1F9tIxAb
4BotGiK/ZydQtRlGQ5UkFnhMb3UjZkRWKRD2ZxEaL6lHoeDSYu6OFw6nEFhNqhey
+sJ0VvLDMx9D4P1ZkXg3g0yQd1AHfHYfNkzzcrje3Rewzq/GHiuHFNn7OYWyeKZq
WeXcjMdsF7Au0jW6v6jJTJHSR6E8KJ+jnJCZrUL90KTDJI/GyTQUWaOxjoBfSQCM
XIm9qdAXEAsjo76iCpRnfzfZLnTV0o5xfqQVmkNOPo8JvnUuWil8W8m3Egl3mWFQ
Sd8v5tjEizb0OXE7zTv6XLoJ+p0RiqBITIgWe53dZRDvtGUaPJvVAI2MeJ2Y/6R3
dSu/tKWWdg4bAEjyq60jerczGqy6RhKvfnHMbWYwwOY7y4Y54lD/e2NCZMCeHKHg
RPp3EeX35LDXqHOF2HWTOJbYZGk2rEN2nbgdU7p87P3Vv17arGaY93YLLTWj0VyD
bBNtyDm0E7Qnm8aGMrlhn+hOUgWxvwMG/JjQtQgi9m5kLOpcSiehAGIqA7k/TUYs
X4XsWlEF2tLXVJpgzf7vEU0rpS8+v1jfF4V98WHWVSu6YNFv1OpP95SJqZlMmo01
HRfSPA1wsVMWs0x4wIrcOm3P/z+y9cYz6G/wIkvN7eYw/tH0PnPoxm4R93CSo9b5
ZL66ujDijkKn+tIn3zoOSLGRD0OHhJPnOHMcqVmC/iYoRStvmgag0xPj1XTXKdaZ
dSRkmJ764j7k7BKHa5SA3AcRY4RzmT9Z6p+V/a5V9OgQCZYvVkD8NcsC11NMaGjg
2xxvfSz97cETUB/DL6ueUngn9oRMTaBS4MfRyxWAH1aJoJaDwsNr5hsnkSzWZmY5
2cbowY5/fy4YwyS+naEamt2KydpBWMtdkrJi4nERzBf7IyylrAduoPyNH6ClrAb/
IYDCquKv5iiL24y0Wz2Qky/0AZ6/USz2yRy/PDVuHrMLkwpOy8bVN+tNJGEf3Upz
BCmFHcS1Xn1SVIebjynw7g5chvgDsPqTumeRxAn+eZESpqmJwUa7Gt55+YaFf0TC
cf35lhvD0p33yorjtSehiffQ0DXVuRWrCFwkzLjxRtbjsKfqUZgUYwt5KHCd8ZsA
yXeQa1qO9kpKz8EoCvzHxXUsc566XJvUOAWd5KFXbcKjRn4YeP2Iy/JMHjnyMnUO
d9oJC6I1neAUNsOGhRDAkZ6g9DW2IxQecmBNh2C/SbAjm7T194Cjv8grOw27LG+1
GOWIFPccYGsp81zuIf2BpCVRFEr08SgGayanL3la5nMUDdM9Bym85RQ89DuiScGG
URNpYhnLyxIZxJnCrFWadV4q5KVHtkbaqZNK+d4JrObdu8KsYW8D8Bx3YNMQ1BZ+
rdoRR4Tfm5fll1YWgWlrrNG57A8j48Aae5dNvVGsufO/BlriIFGyTNNq79mlHnwX
H7HL97BIinvSdjRF0DZjzoXKFSWHjJkZs7HS/RXaPBHf6iSv+uaCJBkotB+O2dVG
oqBJFVxJZLpqcG849fM+hR24Ji8kLvOytZq5GNwr9CVzmd75+7Bw2nZLrF+5yhr4
hpnFTEjqTyyIYMWtnjc9FO4yN9t/IX01Sn5jBP7/g1NVcMCTyfVjDPzCnSux0AOm
hrgAE4ceFYN2P3yzwCa06X1S5QV+Ln5FHkN6ANPJbDNa4WZyHusvdNKfUUEsvbxH
EMNXTUOq9nFsr7NrK8b5Fbo639dpt/zUBnajFxXt0K1NR5i6z6lmP5A107D1KiEL
f0KzmGJdPoGTrQSoOu9YmhRHQH9FV6Gw621iZnqOWYEkURNcaujCVoLyQgrrREqD
C1pQ5aVya4MaZenqfOcvc3IbiU+0dz/IAUcvlIWch51dbsoveN8PfA2Jb1+ahAOF
6mTIetHKExDmzz6dSBljegGnuZDWTC8MLExoNwamyBxUDMxeKoqe4jz3+9y0c38L
mhpacE+CSnaa99yw6TBXKntralHnPswo7hEGzITZhvRdflNDjBJhH3HoaNslZ7Rn
mpOHaSM+FwhueWR4IZhKsn/kdoaHtpBeJua/O7VsCfYfeQQkC+gx6t2lpFbBIbwz
9x4YWkfVcClRWqcBtydpGavvZEM5BJ/YoyhFaD6sEF/Ldl6F8L60yk2KawidVksd
hLzCTJf65QQdo33p8Cf2f7jlehn00uWej6iIu0rsABwHmHVamTjlmeOaNpZANdZe
MMvAJBeRcw4mD3AFdY4HeROT8izZ2dQFnV96y+mibpBuOLaedrD83vGKcauq9Eap
ziiw2IQ+Y3vs5v0DlJ0buoa5iVOHt4yVBDNvufVPpWaqOm5Aa+xVabn88SVTfjDC
lo2YzNUlZx5POo2eCA7glPBfbbKzpYeUyUQv09Rzx2/GlC+9uutbzn5uynyhMLIN
tZIwznbaE/kQHXIiVNQfqcrvMowzljol4EX7szkp8xoPkRZApIeo2z2NgxLfx38f
HyIj7IIbM3nzhNwpi/AVcoxkZeshe5/7fUUgG4Lc3s3rxF3jEYkSMu98z7/U2t2O
5MECH82u0yTPdEo4nehiZlYS8kZFhLjP0mcwZEyQ7ZTy1GuKoiGd0OOJyb8cOxLc
XocVaH96AuwX5aHJYw4eKA2NruA1vxgceS/v3xuc5UdTTyriMkZEWWwZfbODhi02
/GrSCM0Iro9jlHhaflCyn4n3FUwlL+/MUU8LBVn2uf51VB/I2OuhdFYa+niO+8So
16IXO2J6dSwtcJPl2O5MblnYP6Cv81/MgCtuAb04QG6Q7qrP7L0wbTPHSA7Gj96t
wCl7ON40ivD6IzFAWxoZQ+lOHxaExIlWpMd/MxdhbxDChM04aNQW4YAmh/QcvCR3
l+1k/LIr5u8xalnxbGfyU3F7oNCgoVMxUV1YTNAwXRVrNWpkCypzWMhTdGRNQfGO
4fy+VTXL3FLTnYMULvU6nslVB9omrZ235J/eDmkJeEF4fEacZ23vcz3lPjEa0E8F
YYFAwnKswpeBlPfUYFFTo+GdM2A8jCsfHiwNeAakTnhDPdG1qBQBln/zb/NaYY04
qYOkoXxZ4DtiBtc83p2NfzVyIoPo2RNrL9yt4HhxwC/e2cizH3RO5Yb+C45afzAS
kMgIyNhwR/oCvB3MfWb8pB9w/ZIh4apUmVmJzrV69eW/JMWI1P9Ivq3NlG3yUVH9
OjhJMn0ey1rbogMhM2RdAP44EwTTLpzygSrR16F2D2uR9TGlgSzYfRzB2AIe+tHJ
kESsJeEKL5dJsIV3BbwWz4TxTaszgCUj8UXrVKz7bUscUZWPbXSrIdNoI/qag86R
VA5B6yIODZCEkONu4e7Rg2AQmvDXUQc4xkKj/D2+ZvKug7rCOm0Kv4tq/+0vj+EH
0nBWdCakrVCeEzDsutzG1HeGHbwGUjAOKml5K/WNcrsBLz3Mdo6BUzFvBSaqJFIb
O0OhvgYNJ+EFGP/MleSUehhlJX2kNby/Y5W78JeCV1VoCq5TvKPT4V5UIauoeLWw
zdoCuj36Q0QYnVdicAfM/3eHNOWZMi4SGvJ0Y1VKjwgqT9buL53N396IC6zjmsyJ
aReo5/uXtEZgCSL38RiSFkjOwURhhGEd8RlnvKW7YFWXUd5AbKKLWAE9vQBdn5zb
D7SeL4ddcGDyDEM4supYK8nalirklW3IrOnPo/JqD5/itrO+8TmoPZoTQnC6HNAN
zYYYMCvVFRpa/z9lMtWSbpXJcdmRngmO2G3qobBCvjLolC87wXvE6ug4oG3Qf44B
hSR9QOOpVc4x2ClKlu5u87aDg6F8J04HvuKKkF49GsdEx15POu+PYj0jKm8oBVls
7t5LkzvAvAzLMvKkfrekLTiMRKAUwuh+Zb1pQL6Vt0s2XmnketD4czLKveztabDy
x9K6n10QSMY7Sx4x56trSCJEDV+Wr5+0Cxh3N2WnKM2Ot8Xf38zCyh/jwU95LWWn
HAwmE/Noco4xBuqMI5kRaOai+6OHTZWLfh2DatYegmiyKr8E1aa6MTZ3tHfxWgSM
9N1qYyf1HAFdzkg0ZN83IqdRlcnufMhLjrJ3FVXLgqMt4MSZ08yXiXku4ZZMHspj
JYMHgNHQlysuy413AMZTXe14WKnYpWRpFcL+lqVz839sAGfDzRR6ZDKeAAtguMYt
+Iw35j/Cta5IFKVFkTQcaerfoV9ZJ0TKPBQzeq821ztvIPkBeQoDNwycOoPup4BZ
A7YAxRw8KLuIS4NZ3Ec2JAiB3UwEOcpqrXwSW4jKv/EF/+lwjIA/PAWTUAIy5iqf
bBBGP/KBwvA+sSNQD98I+66JgKD8PJRmNg/U26QIf3Ym1Zv90JKms2ooUA7UnpcB
qkn2fCRmjD7yo95KJDa/UoTn8fZqJKyHYar5f9Z98vRRRw8MZ3DwsWPlpNHih4sA
6tnEzqIKKdA7ZbWyoPWkRuHhO/UBeEzfHUc1NVY2JgUEWrjkD3j605AwHw1PbrYe
VGxqIp/EY4nkStO0SlMfoCblhU+4XW6PVDqPqd+XnjLeazGUkj/5gQSyWNKLMSoN
TrKJORJZhRoXIZJdQoycPjFI8rE9i1sA4MlCc1KNnaXFeky8nQ8Ra/BgYsQJ0c0A
b925Bavt3IbRAIOB/qCBacdCDLreKUERCfBZ7je2AN/frYM8BjD7GfhOoot4LXco
lv2U8R23HyrjGV+ET0tBoHunZLpHgOvYNkCQbECS+5HqximQcSR1Vk4NTcIwGboa
0O3fLjs48Q+22oEV/5ut3H12HpkjhzQwkCMSPsQyWnulFFWC84mAFb4EtMNrBXzR
3QPRW/7fcLwJSpXe2w6vZo9QfndD5mdPsvHD7FDdvv4pKS2gdEJkf1Ps+fIfKOh2
iqL6intukfRrzwxn0Sa1n3e17qEq/ue6kJDLdz+FEvoDyJzbMGwrbGbCWmBKetZ/
IuRkiCtLwHJwZSXfKZ4OS4zU2AUyxaVLj6+fO0kxiC5xQR4eFXAwAly+ZUI2C+oe
dlcrIhYBNzHlodhla9PUvzZFtrHcIJwNh/t6PdxbsmiTlkM8hfayY5a+zpHXIHEB
0JR82b+r5kOtCCo+d3vSbG3MsBBGj4V5KHIfMoX4Xn4aPmQiPGAc+HJ18DUbxNKD
CR4LXG0QArJFkyHs4YI0hp0lS3P+rj+Eo+efd61gUlbqx0M0uYaSK8bv6sjOkcBa
Dv7fFgz49tn3rGKu/Yx5u28D1TcGrpo16OIrjoMnYzD2o1Vv3ynXtpAZrGK0x5EG
SpvKBIgkc8a7+2UGy9lmZheUm/dr007ZaILR6sKUTmGMDcxlYSEuTWoSauymrMsd
yZeFfW/4jnsHAfll7ldDu/FC16MfsF8yc6cr3mDX0SpugCkw/ShQh/PsKuP77Edf
7EKx9bBjRhIVyR7ipRlO7T7hmXz7sKDccNiE6G6WIKm4/k+GE0YomuVt/XkbMRbs
6KfI/Lz0ZJ4lVss7qrnqYXM78O5jowb/RYo2UE11XNUWMy+GUcckfnb9MXszirLc
NnDe9BLnj0ZtONdYUqFUD5yXFMmCL0+xURonEX2wiT/KmJDcRdbG+Xhce/ecsVv7
EDnliBExnb/PX/GpXqd19IQ/onyeruLWPPkPJpWFwnGuoJ+diLNc5MrZV4kxrpEo
psAaU7BIQAOvDUgBVJND0ijrOBfU3VH9w7N2ynQNvAs/30vzAz8LVKh2ayMUZ3uq
M5PRnIAccaUrssg0iJJ3UYB6WHcHAC24wEMHagMY7Eg6fns2ZsddAV8XQfiF3kJA
rO9nDuhJNhmX0g6FvVcrNjXyjP0I3KxfplZb25dyZ1LbtWDSkZ49yLn3o0EqTqQY
Fws4iQydeN2uk1ues8qml0VdlgjHpP8S1MGmSTjqgFCJv2vtYduS6dAobNH3bLjv
O272G/flbLMCnz7XOf9sGJa3TIUrAMatWNzRVb99gbRsVEy+qIjcNdYncY/wdotl
A3QMsgnFLFs2oZyuTIAz75ifOyxuTzbAlN/ZPExy7JWztmCX4nHUfB6UYohJHU7X
VxuCrTEdR/h8tgvgmYrGQem1xrP2Qz/2Xm3viDAkxtLZWcr+ag/5GGt5lo3Cu4rq
1G8Lkhkuk/psgCLJFmkf3ta+MLyUXKuX6IMAkoJnBgBZZjgbdkw7W7i5W6uC46Tx
r9BWaVEJ3syxcYsKo3XhN0dLeBmTH4k8FfV3F+lnVch55g93NGuJ8WT7EwiRs5Ww
5Pkuohw6doYWd0TceHmm4UjSH2ehJbyunPOtewryjnYCDxHoSJj0P/LLAFRYp+AS
B2xV7SPtlMwe0KQZ30epqajogRjb2lypWUnJOzlNWzAdUFmABkVia+vAKA8ta6Fk
ZX1l+2LDUfoXNuuHBIXN7vopgRhhxRBusLFQboXxmS+dECg+Ia6qDs8urHKWOmk0
CrY+vQvU/4V0HNY+HCbg43NJU50q1esNepy6ykamgflg3/Vka+uLIPNxFSJAaJGi
ELE54ZR/OONEtv/I0oNE9QmOu1xAi4KF49OJBB5vXSqvUIqvf33z0JZGVMWgTdkz
3Rs4K5WXnom9Wd34FlkY05gv+OQyLCe6ogQXIPktyzKMmuYlExJkhV4GZIDyu3nH
XUtf3zm5zQtQt1IGn9ru2HLq7ifybzokxJ5bNEQvgIka06rEVlDNvh+d/TmsAIex
v/fZZY5WJeQZDiIBXwLPAIah+OUENzVIJ5DtIBYcjBDiSBDa7QpS0OVGSmdQvpNq
pd4ylByJuOSjZHuh0A7B/MEGY2hdQwuJ2HzL9EX8yAvOcZQ6L5XvnpdVf8mSmKEk
a7P4z0KExuU+cLdgmKa0XGnITe/+9PYUmY0eT6fD9Y1mNiUduhpbbT9o6B/aBkU0
DGsqi33yATjSUv4UW57YFq2STbvv0pTWNlZNEoyV68KpJ10tGql35TMqur1WwHD+
QjmaapUt3tdzq9HpTLs9fyEIx2rH2KJTow4qPgRzt1qL44lgQeoexvV1VNDNMVWY
IXjw+cu/DlC5sWt/nL2j7CDX0PHEb9tlf538ZmBVCDszzArMVV33BSGniL5jxx5U
VGakPWPiUvnj96quMiVbff+qYupk0xmGPRJo1W49vchyKg70cJoNjR66j36l9EBD
Q3FRQlor/3kFh3/FcPrrxqz4/yaWvadf3v1k6W1/iRWSFtjGchFoXB/dvSDZC1ID
BRSJ6g3EMFfJDPP2/YP/LFkoQ0t6QR0RsvTHx3GKDIo/J2NUiAhfMEfeYMnLpDkX
yIZnbLL171kB3G1TcU3VF6rX9TcOvbNEKWGaGotbmthzjmmdXOMp0tfPOtXXAytE
Xrs7OMOa3PElp72pszfxosYfHkjqeqhZ7XdhHbnFEMYIpiWMjcMPmzVhEsuAKykB
f/1ggOptJbEqO45O9DDQZTXwFu977muOOq4/6k8rBUD6wTr+fLQHunKqPSRoc6iI
Ybe6Gp7Ek+30h+udSfwAiswHpXA5Yz1p8RJ5yaqC5ZU/sRCuz3vvYo86UM6kvcgR
qO5Ufbb78+5Fw+BnYSb/LtkmlZwuk9nWfnDuQSl1h3YcFIzeXuLurlVGSgE5EUXM
Q075ZFYtk4hpwB5mSLEIg5HJJOq3Su+XjB1Tj7M68sh1h1/QKgmxgS31qod7DKPK
jgRy93z7iXS/pgcCXFXjai8QxItSSCvHVkjPZerv+OpTWh1SxDeWwJpUx7+T9QiO
R7KqJCh/hJM9IOvYoClKr603fYkqSZ9kDIg3Ye53fuHqdv08+BRZJQkLOHr6Iw9p
GitTGZrhTS79Z75Tae7MyZdJPYtipTKMYMJaObql7aHpPa/kE2OzlMmrG8ulkMhp
UFfhW0reM/MSmWK8qAP2mD4iH6NKPlgJrtnf7gxmENMdZeVgSFxOkaaXamh4hfzq
rNyLd5nG1igUrO4K56AE7aqZwLPaoQQZh/WmGNnaqRJLJJaU/RTVZ/03JsfkwckA
WZjleqa12+2L4630nWT51+U0pPs6SdUbAabdHh4HsCAowymNj5msz6Y3sZoaAtJn
BOHHC9vD71DRFJY6xL4K2Z0X43Hgf/zk60ck6WHGGxMZF8NAWvDoxMRP+dn4fuFO
LMaaVvPELv0NmYw9f89mwTLOnlU3JzoUaZ9n3JCaoT6O/kH7WS/MaIaV/zTKu0+6
P8i0fCOsMMKpRpqVAQ7tawMkYmZTaaJWnjJXwr21eExOd9mIcq+CT4xaeMAqn4qF
bOAHf+ImKxYzmj6cycXsrX1lnU4YMnmhKkZggaSz8dpkPp1+QlIJLO0j0BzOV8oO
IgEbeGeKVg9JMlxeOiCE7dB+7z9h+fkDDQNzRhaQsDnIHwRyuc7hbv82yMlteYvD
itXs61MHIcRKWW+Js21Mz2rrqIW8+hu7mQElLxWUKtkI6wqJggrPCa4O/0F7cJXU
oZs89yKOjvFNllN39v+c9QbmF7nidp7CEe8/LwyAuBh7dd0gNQjfvo7lNnmdb8QB
818SPRNfGQODsQUePoUKVkZa0tzSp32IyYQ/U/87/yNEU4C3Vk2VDIdJezKYCQOj
GsL8LO7crT8bD460CEjdqCf/Yax5jlpBm0jYMb2cX7urSlQZud+e1XFm0OpgXTn7
TEXamIMHhVAPTvmagfxfn2svgq/zT4TIe35DRUnj4E0h7qjR7FkqFxTbo0BrHpue
jjfc+SwfNSIq0IT6AX+Z2+vX9zAg42EYi6mkx0d/R2/wimgbXe9M/6CENgcG6ada
k2X9nOWZYxmQvRBEteFehvHWMXw8P1FSZWVA4HdzxQqJt1h0cfOENQHc2Dp46kQ6
uLfOIWQXDGZSEO9QtYUmf6p2nmKXY91Cg4SvGfa8dHnMTaYy0ugSadUqNZaIxMtm
VSgkC/NphxOccKhxnNJJiWy4DQelAxRWTpKz9WgLICht+9j2llcweOfd2K31aVaU
IfX9V77YQCSstctdB85D80jNC/t5MKlKCAe/ka805oh/ePFqc1f+gSacRcg5SqiM
I/8+/AQ94llhcGJIUmo8WyUVQ4wYzQiEi5r3PGJwTCBbS/SUEF7vZMFbEX1hzyKU
xCZQaV9p4fTStI3HId9/j16rOPt2KTCUzJKLkcy/JYxxrx9nYt7MGdlIddFe5v8z
TEnKF6wMaY6x2dBSm3+GY8MMaU4ZhYxJ4+4607ge80dk6D4D8ZAmUZiRlsk2SLqj
ZK46jJhGlqJxlsAzp9sUETkAWRZ43cPiHZKzBNastnO3/nfLBL2dhF9V5JmvMLZ2
4qz+qTdEHHYoVULNJy5kMnxmtzy4YstjnTEZI2z9xmPp//pSktUB6v2WpWkj79ZJ
NsMh7IgrvFh+jBBwoG7JyGpS+LrGNbYA7dqGW0AL2Bra4dsR3ylV2HulDMxz96wF
w8+IDu1A6l1JsxLN0oXjryXi3qe7kda6zcaM9SWkFFDiLVvTuI/UCaEl5mnkHKW4
RYDzoXfXIaaXLRyrkmbd1C5SYJDsMK+9fllfczNbrw6euaeGe/eTPzOca3m++0sm
nLiYuGZ3lXOo4AU4pfP1/GuB/sfvF73vgzlmW/J+SxiG21+XdPOdbVgVm7EJj+K7
U5ELg3Pq65ijwqkQGJy8k+Gvoca4RaGizICfohbMFQzZaUAF2ug813GB3PNJc/+f
Un+8RoGZAkzpjKwPH1geCJKJrLJjjl8zedqw6TlkPOAjZ5Zw2fCIhWikx2+gfNQ1
RvqFR323Tk2WfKRobdYqeyAmxzEm3IDNNP0F0n9tXmjU8ikM/7QeYd30rqWwMhim
5ERC0i9Sg/aqa6xaY9up4a5f3AKprXzlvKmPwiWkQauPjb69cF6A1g35fuIRECzg
PM0lUUQGNnYjPuEwm4QIG4pg38Ar2FSUaZFAGaF+EqJd8WG7V9Amcfknu01rm9KF
OZfS06Q8Um/rOW0z108H/+yFwo1eAYqGeZ2xKkF0xjG5cYtdt4aVVCHoO5zS7iLX
hQPk6e594FkCRZ6tjTj/lf8ng0z9jxOgbDX7g6BAows3coRpGWPanSgv/CdDSkgu
9v/KxoIM4EFCJblhKnz3zckiyaSsV0VFsHqN9el/vjybwBYbiXUM8xW1sbJv9waY
1E1jH6nS9bJg+TGnC2ZKjiPdX0i0PFdabNUdrpoOHXN7IEI52n0vwVywNELtv6sV
3Pp4HInKF6YMI+bMmUavV9KDaTcSuks3tkh+mTl/bNjoLN1cb003h3KhOSHnbSXo
qAx3hV6hXD16xQAa9VeHwCuq4KqVcxyfeex1q1Pavu+jqylibiVc8/Qi0CBQeIvY
zssGSCvvIZp14Zn7P3h42r4NRc0buTZfewk+FDN+ZAS87v0q8Vubmpxz5OgcQZoc
ijbH1XLZoTO7CHCYNXIp0kmPvxKKk1R1i3gfWmA4VJgheNyIXtVJnzR4iT+5l3FP
n+TcGXD0xXFKLjJWBOs2siumV9Rsis9aTGGwzLtSJuuLDE4WTCGgOfvGXuo1uWSE
1tpe2BFSYq/9ln58YPOSxxF+LMCHyZRd1DgDUojBuHit7GjP4DtWfcDbk4RLedtU
DJ0lHqKxIWEKjnH/b7BN/vQA9wNp2mZ9nJ4J+lpqHIUpdebzbveFYl11SEFdUKHT
B/dDmuPwoQCer+JWKMmjoml1heRlt4YtGqBU7m7bR4A8HXRNjE40ef9n0OzbQ16c
W6t0RdvJb/qG1cRZvVto9vH+HNteWbdXzhshb8cKedsjQ1LTPTL0GiyEFzqfV1Bu
Y1z6tFRhW9KUDkYLgVtfmfkXk+bRyszXLNoSl5laCPc7ndy+sycAOg6dAkKAv2Hq
LGZYVYA5gnjaLIx7VAAcfD4aMGRyyH2IXgqNJKQfx+l+wl8C2qyRiEGEv9Ntb2ej
UkTp5TeZv6Uxf2zJ7m5xZLT7oApn/MokbVfUiBnyUUAIK4oZdZ5z/+WeKiGLquux
Pyyd160GuJNa/cNOCZn3not2scJcZbXg0Twcjp03QSiiKIV1OTB+j5SCDj4N9F42
Xr7M8aszDNMNQuOr1m5bjdVbyVKuRPAB5oFkYsxhf2gKXbzP9USYB4GLQfWVlqbL
AKtiYQ/76gJ3DID2bswJGIXOURl4nGqlIIfC3sie0RJLTkC2/h7E0dL1KRFbC7ip
viNkpcXAyDOqcaelQwNVgq/qgfIoFpjZrPjVBuCJMWwoqWv4SwwMoRcRwejfxAkh
rvftKt+iW3ommcS3wvbl5L2xHODUoi1Kemj0EGILbkr19ZmKVCekAe353PFHi9Hp
oBEqZTTpgFgL37c/UbeermwdUcJLqQ6sVzkSTf7b4rRn4SskcPjUJKPDXe2HZgSu
EqQe82ay6Fgmg9rGOTRvj3p6LIkxVD2pq85cgS+YwOOGF4Y6F8Gewbec6SY1PqmF
h6/BGU+jgNAFpU4pzGNvV50q7kY/AfCvaEY1n1Qmh3j1py4xT861tojFKVueo+uk
eJgRkrF/4DjnorodYpAQA/4wr9z81tU8Z4QbGPrux4bYSADQTRBCEwEEluzUEEro
DjaYvOc65mf0QmClCcQuVBBzHdy+XdD37SHlQL+tNo48PDkmf7GzCBMsRZ2NwmDQ
vPDIrCWD3iN71Yk0nIkfc7eJUD7KmTPGnk6g65bD6w3fFyfcfmpowKA7Yv4Xpa4i
R3Rnj95YAyRvvR95TqadFNdgx4K3DzANUugIgp4kxCUq6RGaoNbuadNwjqyTntox
jiAF/mUo1gn7FDSKm4mwKZ/8i7WyAIW1XMkhv1R3z02aewWjg3CmXcE/N3ll6PL3
sIlTugZLAcU3mIt8zkvw7Xh8fHtqeAXY6uqmb7YoaWKUflTchSuzoJNV/XJgTu50
pVexLnYjMezFvQrOqAJ5RejDcsynSfO33iRWRNa5PEFpNFU/ROxboJ2KUfnJEkKR
C5V3p+fqP36Z1Y72Y/rFEIr8H+mHSh7BDT1xEcaZuhsdSHBhhCc8egmGs6pQkZDz
4KTiL4MsmBoYbMGPrOLcRq6kFd/acS741ooIkUkEmhyuE9WZ4/wT02o4k0SGxo+t
HxtK3K1Yv6GV3vhiKhdKYKR24EK5xxJKCNeKsgriQ7uL0gZan9Jiok1YZRsWRXKO
jvVJvFPJC1RD9mx77NuIEkMgBcY9sakvvjkjEgkiShIH9pdiCQCt+aXc6PQJ5HYa
r0LAt+gVTNX7neXZofOnO3tRL9pssUYIWrbFRNN56AcxHjslv8qVk6JeyognMU7p
gzjwq2bi0G2ViakP4v7/R+3Lj2HUAo35srBZh344cSS59ZN4nXUpIb7t8ZQwzW6+
ar5Vf+PV73NNQUtM3G9po6i5KWCnqY30jttAYi/YD+tupEelyavf4ztwqOT47w+Y
34QZeobcG88C7waTKZ+f7K+gc5wXR1cvaFmaLzRjfA3pP79oPkdt9vM7rEDNi4kN
qql4FFGpQW69zZbgHPM8vYssg5Xj5DrCiNrk8EPc/L8NAHPe8+ofkdRZ5YGqRiES
qbfEV6eBIi1TV5ewWcB95GCnK8tsE8T5KVAiawDt9cw49a8fX1Vvjxe2Grjl8ySm
rn+PM5OOrcw0qeeaa5hhU0N0qwJ17HPsud9t6IUGocwxxjtOGhSdmEXAAgDSIh8I
XHSZldvTS2BKnv8H7nJdTWl6Aju+pVytZn09SU+D2ASkbh2eDO8brEryctCnhyo1
a5OolnrmrePLxgbj5XkStzioVGLQU26yBsRa9Q65KyQRCu0aHMk3PaW0PNlZ6Jfd
qiLXY+d3CC/wmul/32BroHFfYeN63K0ZUd1dSyTnkYb0KI+/E4uoENu1Kuku2qYZ
MRzSpVd5KdkpiJWHQT2Y4IpXCtGs7+ZmciduBwMTP3QRr4c+9HmokE5h77whLuT/
05w68aHtZMcIZfN9ujUHsJbXEpAumAejw+QHQxQAvzDeQXk3vVnAftvjRiByU0Td
+kja9A9aDv454k5oiNjYpDrE6AfGPGfNIImeG26fJ7qWK019OuGhSe2K8BM5ixIa
D5E3mYEixyQqeQqe5Pzviwoe9mb6C1BTrYMYRE4dxz+kqIsrp8nTyEZmc/8QQORY
59MAeRcEiMX3Q/ne3+0cSFDalGDxLLQ8QSimu+LnIe7u6ql3y7b0d7zJIGIgVy0q
8bpY8HhbMXqYyVzf2uS6iikcEJuNzLLbxAwWu5eTKcax5VLH9tUcy3Szr5Fnkw6/
adL6MQF9MdrZyR7qBdhaXPhQ0PZYfRyEp7J/GMgT4adP/doZT1EaaNGmGF9tnk83
IBpTpzGt17WAFjOtvzoJBqLhfVuHF+3sJ3a668WL0zypao2Vj65mWY24BRxuQNty
9QJRrjjCbb4ISVTEGniYW/VeVROSthikHD61jaIf/yDOmITdllgs3qN+2gFVog4P
3KQ8bWp2ml8plXWXj4PV/KBmlKA87LxU574UTF8WAjpr/5CEqydJSKD7W9fyKIFw
mMJAMAz9djeW/voOg2vXlZSmfjQKsJbVFo+//vBeCyOE5AyYGcH6aT7xCWjqe/rB
mU8Q5j0wa1bTNIMMSYBgFlP3ThjK2FAr07/fXneLmHvqE+RnM/XeiJ2++45ezE4p
4EanFjWN8RRflRkRwWDLNSqH+1c+rnelDurFruJQqy/MRgSzuQQgZFhG2X+CYoIk
ya7m0WYwWMg82b79jbbwtBXn8TehKNmPJKAF3nRQNM7w4z9vGGhIm/DPce5Mm/4a
rE9NsEfMpYNGC3jwblCrPk7ktw5vWY9w6rFuZZnP/uW0ieHNnAmt1eKwOscfDhKB
gpKpwuL81V/BcyVf91h4T1QayBk7750GeIwmcXvGKcCEbvn2M545liSE3eUXSDZS
fLy9SzS273cJtr5VNUaU3KkFCaqut7Uzn1D7VYu/WSP7qZxGk4tHGXYO19o0W4P/
lENb+kVQsRmMGCZsqdOr5KILS4+k4m4w4ZYg/erPUQ1NiKJrtF+1bQa3SRchIZ4q
BrkCiFhC5w76JXnyTn5ELColu5raSr3AafsY1cV15GtQELQZ0GGgB4XYBJeRCUTD
asUn5noyYYFpFUuwSLBYll/j9bIhDw9LfFE7B+PtOSvXabTiwmIUvRz4wtpifCIR
rGDP5bK3dgbUwUg9OcjdiFrbTCF8hd2Pk4/UzUWz1uJ0Ybrr2PIHJIg+MBCc7cre
h35SYSngIy+W1T2arsdvFsDaViVMgWvZPjn6CxEcGP81MoLyuHP5xIG/KBHX3yPB
pKFRQfteHi2E+Yb27uFmpaQoCviT4p5DEEYT3o+sHDY0U7/7QWYyXRoZSx0uKMKu
1duzWdjOl2FpoKrbUvrcylSeVTA67jhDPautdIOKowJd+du2RXoCMqttSPHPaQZE
zS6HA8RnlrLPZHlMKYoOnDI+CpmJQNZ1WmhzWF3x4RePDfqSKWMMhRiGw0WEpZO+
bm9+FeSFjTPt2Mj/yLDKDn0lN8FiijPWH51+NO6EAUn1nt+wIsEIRfahg1hfEUzx
9/u3s2wjYm7vc7JU5DKv7dSwQCFl3nehZ06Fq4XtifItcMn8RrDGVovD383ochUP
0fwlpyB8TN6yipTWW4jsoYKZ6w9V1tqIpljmMXm4gJxDCEITqtJkX7V/KXbgHjbg
t4uXAdkHf/JOtBlqWkiyMW80GCPgFuZJYcuErjZcXQG1XGf21+Ptu1RM6XAk8WzN
UnhAbNSo3rhWDRLt4vNLbOrPuJpCihmZv8ktApMtwnxO1pxBNOxN/uuQYj0uV172
4l12q9Ll7M7pNWEGIDY8XjpRM+h0GzLzhZBYo8i3Wj7EidMTqZ0aW7wNXLJ65erw
E9bnBuQDpnjCGSPEoSvYnbEUoQY6nChq1SvbYkxjWaMg0vscPUSvEBc0+qVHZ5t6
zlQGFZS8k5r9FSVtfm8WdL4XTDthR2E+WsGFLkY5pgECsqv0K6mOp+LuR7RGsbxd
0/cK/e5EYix2/GGY0HuTuExhLgFPCyyOKepVEjLNNmA2jm9dig/DaMJT3BlMK80f
l47lvJJWlnAdWm2HR86/O84tQzT4Vn180v3YM+AbIDa/sxCaRd3lRkvsJyReMVds
KivnzrejWIQSuCwOKgpBOVugZ2vqpgFmtD2UTrc8Vp0JWjxbrX7akdM31Pj0zqms
RelFO1FXvGTJg/F/wTBtpWcvjgpSAadwy/irT2h2XRm0wgazc6bChilSn8Jno7tu
vVSaBlWN2Tm2DiMbGfkXdDhuxROaT5oCA84cpkC+Pq1LE8BfQQlOPDcLS9HbFXxf
spLP4uCab0ThynueTOYKl9/5US8lwvypPeFYGhXGPRnsCmP4/T22OQmoiK0/vcnm
E0QVvXT0Kpz52aCViJTnNAOdgHH/ulKsL33XlHUah7QhU+95PKKvIM/M7mTg9FCx
UHvkByfRrVQDxmDoFjRo27AglZJHAIYdX+87KEfN3jE0TjE2QNW4VrHLZwg9BD0S
7iYo4XFCLEIDYQpwVzBfZ52QL8GcoNgrgWstzPsp8gCdyOAydm/4z0jed3AaShV1
gi4PU8H92sf4TPbW7Rar1Pmb2ob2Fjs/QLSmLmThh8SQqHpg11/3OIjC2HQZrZZq
RPOCKN985w9YWcKhFpnCF3SrfwICLIm3ZaGUqmdZGctBnwHMjxRVVLrjGtbEkBxu
nZ51tt8N0+qT8hpeTuU+GVgZWkz+/EONZzMrMHXYI3rp0eAT5JAh48Qv8xTl+MsD
xAFlCLTfNrlAkDmvhON7quE+bTNC/VRskP0hlAsYmOxTXu0LzyNlH1cGKTAWvofi
mjXLiCWPws8/YzmBHVgpURrjlLLSSrV9pPTc33hEkALCpVaKupKLN0rFuCLqw4mp
WJuz9qHmIl1TTckS5L0zLWkRiFSwa6Gz2kBV54o4h7nBvWJdQ7mEWxMIMKOvAz8X
qWRGjLF4tXWNSoWFYtFHUO5ZfPkDbr5OExzsrgsTgLUL+nnhzOUj5H+Xb2a0hqYk
s1f17LOrusha2sWOIL8jqTXHTqEVA0CH2Vh3BDIU9OEzF03z1lAwYrWtviTRGbMi
sFlhhKD87lWIk5cGByeHm3oT2mEe8a0ZB9aKAyCAnjJ4P2+1Jo0fWUFH/dRY7j0w
hjuQbtWTtbkjc0Te1nJbnZYnZGfp0l3+F+FNJ6t0HUACrD4OBXgrZ4LlqRXl+73u
koUpXRe/JOivEQIl+4r/W/+9Jslm8LqMSfPDGJ5BvR7Q8N5TtZmOuKpmwp9VmV1i
psoDbEExjSkKaxA6mbS5mD2IKA2/0aGoa5XHEkNK/cF5mmSGzUucqD9uVKlKuAHB
8PBRfhJvFUywplu8y3UfvIMOMcTvoP+xle9A7QgBp+uQIEZWM9R18r9qpk0aD+OF
mBeYnobRZgtejVlZWlQQewvhiXLhVruupjtaiBBKIPG+n0gGXwkcx/ztOK3RLn6X
4DQzFGQbiBqql8eX2npALH6/kEk3ZxJnKIXTXd4xkVllL0SjUndNujv9BgHigPbC
Ai9X/rod/K9DumGHZPun/uuzH/nQI9VZRM4QhR7fppwvxcxkbxO8BPjlttAPcwQh
qOnn+GOisP3XJvAqifTkAMTQainjKCsv0bTbAVo5W5X9tMxzygB5QOL6/ZGjJAUH
+eazj5wIBQzeN6LJHJAcKdUB2mEZZ8nLpMLBFn4+DEbQDYdBQF+BKSg3a3ISYO2/
QbpksGNfb5NSmB/m4wxtz1zI8otp9rqIUqKMfD1J8mEW8LaFZFWJWb/8Q8SO84Sc
4N1+vKuYQZcGmX0+Rc3+y5p/sDTaHh7jyvxBOerbn2D9Qj5VNcVTIizA/Fys2sv2
z8FqCakQRnnSVp7J3e/OWPsVFAes88e6WzU6Wu3bGhfJ7xKfCm42I5MTVXS5N3UJ
69xxgiDaXGmq9H+1DB/JKvAYvStqsv+4UYobf18bNRfM6bHQNU9CXCcyQH/g+BCf
SvB8dUkS+jHv9b5diRm06ZVDZhosUAciRTBasoZBLUEM6GDBEF890RTDLAHBqgq0
eYCgyGOzpbaiJmwALyspilxdqjK5Cw4xlb1asB4AA7HfMcAWSGxpmt9RRpN+zCDC
xWDWmb4Ep++pH5ffc2u60Ix3D3UugxCmKGFua/Hqxb4n3qMITtFmMHITYrAg9dQA
rCvJa0dNk3pZn3LEIQwc3CGnn8WYk34B1a3j/snBpAa+hirjYOKflUxwWlzYw2nw
Jkpgn3ZkFNn8aV+2H7+0/559hyIzFy2AHaKLwF+VGQPL2ynaZIiZhxjaMNZi+vGh
Auq7T/G7xqrY8t8+irXrMkcwGT3FaXInB3ZFXVf4MKud3xp6s1t/BB1Md8+AHwXp
E3FFwWtmp5c1BIiUBlAKShF5tZ1UnqKm8++x9dYqcFhTIzELtM7x0a728YTKQaLM
qnvoigBIyaAL0XOeEeEsRbcCqCDz1kATZDAcH3pdeC0nBy2wwc/e3Gblb73wG97k
3QVnUky5tcHP5dQg6O3xrkLURCB0U4ASuj2pYxnBtZKhcFJ5lOEhGnYS+q05gCht
D6/h+TytAKsOWJ29uD/v173KIIsBbRLOZvDZXMqEw5tEsXnBz4pfzoW+9RR0Tpwa
/3QTkG+l0WXHzvnsuVjcbu5apab2kN6PXCH5Rlaem7wUgTMSXEE2ceuagwsBP89P
YaSpHRgO/UPuG5mB+UA6dFiFu66RcPpIgPlew/tExUtLe5Zc0L+Xw13uw3VP3/AQ
rEGQnJp5Th0G0wJjeamuWxrR0ul5Fq59NGdT/O8yJ/qsW0kFTAfvLys2uuQDZGtJ
3n8fxFx32EzOwIcyzq/2qZD81RTE5tC/0GCd+QT9laGCMWMX8AZMBZgRaGNLxaIe
2EO8FSbuiNUqtQ6vUo8k7LLhe+57fNwdUIZ2RUZU35ilStZrrTYf0uMpyl8DU/Hg
oYczAKqCS/WRei/blyJ/HXaHVp8SZsEDinWXd1nDNGDo8oD6JowWCBhFBpDcJR/Q
7jOUWn23cnra4jJ/59b/7CsP7TFmjNgNMXGQMOea/5xHYXhyw6ioAahvsenpbrrf
okBToBRDBWQzRkPody5DPeNXyTr5Ck7CU1BIcsH8ALIlWqllgzXgsU3E0CZgnBxF
Ap4w3Xwhn0vBYpKnQvjoI7DQLrrjpWRFdnUdrpf4owBcBmczDJq/k8G11k8QIoxi
HNU7ZeIP9p+B0C6x2kTm94OWFh/lU/2kMeOg0Ep6FfSFgBgZwnVKlbXUqI+tcJ+Y
xuf5ejxt2AIJwSxn8G/EPXjDBi6KNB0lP9vpbZd0x20ArwdCsEkmutbLC0ToJe3D
Au0C0EpSAgTpeOkYvOnZG44HbueMZkfi4HQuXmzhcZZNVqEaDwFPwKdACgwE7IAz
jiPQP13lujjmzVTXK/Zon/XjXAbGOuRR3aEQc7k/A/9VWX8EYGjp64rfyCfgF0fq
mWBtgVqPXWwKHCB1SppvF6yhzAqMf+chSfNa0ljm6en0QdkY2Vlr/Q26lsG8Iiqv
ankBHXKgrmHfXEFbJRQCQtYzy+g6UP5yq+hbiuIiIaW1/h98dAgtEd35FQMJQRyt
uxGBvupzHUaYaBfUMOmWO4KWrpJSOmAiPhyU9nQdM2/HG14Fq23Pg8g5OwumPt7r
n+ER3qd15j2uphB6Ngl2zJ+frd3U0dPSD3KZ2RZ4zzyOyNcYmYOTcNvkBH5O57Hn
Suf7Gn3FFKdF9UfR9oSNNJPpyZsNGU/rtqfWFsCXSJXaQg/uVrxsn6O9si1eI/67
O70dUvOFNqNwAgtWp6cSxnAH891wCmqbu/Mns3evTMhd45jqNsZvLqRvOmofgUcz
Z3ZkXck0PUoiRVk78qEsJJxIkIDC4AtJkgzMNR8Ib4B9941IM8Gt65pmRjHCaj+V
+w2vB185K+14I/PQqYGSkR/PBxebSkDybs0y/eErsPb86KVaHNlSUJvUs9J5F6US
rm7iHndz53TMeUfu/aaUFIlq8NKu0Rlz/bXhmEoZ1zBKd4179e8aZnv3M5kt6LS9
RtqQKHfKuxgWi1z05fMj49SjxhoBdqBOhoCXwITrcnSMeE1ojjGaPYo2xXtVJOxG
I4V7iqDg03fxqKRbxvRUTAfgsRTstSU/Kz/twCORMyXwbZWRrulKFcVbuK9WXRN7
yVdXoDi8m21TM7wjp9OeOI6eKwaKrT1Vx55vM32sT+VdK/QASqS/sDSMS2y2C3Vw
c0XfZ5JCgkbjdHpqJpeBiS9ycLuUvSxJfNTn7juCVvWyugyCd0ocGk7F0YIwLeWA
JLD8APAxVFoVjGcsXJDYJB1X9AGcS9aXHaWf7gJ9dP1w1XK0RsH7jLnsGiku8TWt
bIMNT7i1VlssIlUXMi6/eyFKacx6hUtZz1M1dKnaui/mmut8nBrYcxHITCAUoiex
2nh2l7o6wajDDsshiX/uU86UPOfvj9qYEANpl4HGEl7U+in1vSReCmZTrkx4AXtw
k6/b0CuWIfzXIsvlIGFkRgCyD2eVjus0SUFRayBFOCSRB9rzyshn9QUxAcO+KXlp
Wr64hSM7aIEHAid+9rsAJHIyelDAie9mVImv5dunqtQ+imEG8zaqS4cZkLSCUauq
/z7R2uNXSZ/keQB4yKzhaE1WBVcu+uZET0AF/JYjh1xMnWtjQz6wjRD2EuDaCYJo
qk5OIcg+waNlJMuFpHy1C38b7WYiyGhjz7ITBJdlzs7RsjYXsXMtuadMZNsQ7p1K
T2z+vRqRtZwIWN2BpzlD+nWt9EC6aPLdDhxG1/16oX55tASTxr61HvOyguk8F9g3
qbkjCQ7reV54yqDAuiUU0+e99YmvtHzlXOG1Gqd1OEHmd521XZSwhLirGmTb+R/B
fylWoTG8Pf4FNOGb0oIe5LlKGM2vNsgy0pAhNhhZH4faDWhoR45t2ZggWkWzSwfo
qEzgEMGcEZLP5xYqDay46M4uCOjgebtAHNvVQizZpX2asvx1M475sB/J4EfvsZU/
mM7a3AZvpwJU4e0NkcKPgqnS/oz8xE5Iywd34jzUA/8qp+C3CNE//ZYKkRMd7a67
BmYkySdPjjtzyERpcewDC5MQjSShUQukfHUmW9aoH95pHtrlwVFqRHCng1RfdOmP
DEUrxIQow20Ciidf2KiWEUUIOsZ75OFECdL2Lfr+9e/ohJCHqlr6cOXr9YOJxFk5
A3lSDIbgkNXW0uE79DWqUPlo15suTOj/GDfoepSugYIoI0vw2HsUmCdkE1X33zct
0R1RyzCZYwRP510ds7P8PvKLvN+nRfx+mAUgjCWUKDByxPUWgj+gpcxtCcStTZan
ym9FSPmkO9yhxJrRYHAqg3zwbR8yIwrb1T4FoLE+4JTqfqKI245TzScXYsANG7yo
r77PUi8oNN3r0ujsZKQUVN8F+A8tQNZN5UMQj01vPIfTfaklJzDb43zvD8Us7Mah
zyYaT/sALXSWliBZnSDTWlVQIr97pSxZ/Yx8OHbYcaD6e34GVtRTr0d6UNsThONW
XtFUdVBVooDL97Jd7tzBvIb/UdZuucNyMUOjlWP1XC9oxL4IOS5WNsqo5worDMjw
Ms+ihtds0gmZViWjWLaQ4xxIRspyrCY9DcpApe6htfCxZB+Gp2/U0WA6+M8ysfm2
YM40oWjoDiVGQP5x4i2Vp8Xs2s1s6sq9QHYITLJHt3+yI73FvOW7ATOHEnJ7lpxh
mehnBET+Jhnn6gQ479rdqIWmhCJjtaIk35TKquMt5SVbpuKlSBU4RPbTn98bJBj3
ByMLPAfauScq+U3vVvAUEqKb591yzhcQM3GcNPMNq6j3ukztOX8np6tJGhmczPjP
p7fA+scs7aAUEXxJZMJc5rc8s+YWTRKwY6S26jtHGhfXdveGUtOXyf9nSp6RjA78
BJF3W7fZK+imX6Cb+B6AHOe82yPdmjAKMvb+xliYDyt8bmmXPete6hR0E7WoM7WT
BYT49co/y0gDAOkcbwDNCWPFP09IQp7OTtrCUV7SO13Jovobuvtj1Ty85m7AwBoT
xMnV5bVqBJYRt8HGdvML+j9IcPiilMoEpbtCgUgkCXsRR/p9EvW/ThCDGSpgDmG0
H1fOH5SVi3/Qm1FueQoxXplTU3/FbdA2D0knhrspK/BXCIZz+ZoEXKMwQXJI8oNm
bX2W0SAycaYmIKc74zTIwi5Bkw4RxJeBoLe+964dzb+/2sPlj+qpL+mQe00NyIYt
8L7/dt2qTbLKb57SKX/7Ly4YIeCNFx2qKpNUwTTKH8QfH980ZSblJnAvylJPat5e
B1xyVw92V9p8onGc91UJVJQFuL0/WdMLSQZzw+koR0F4OZCpJtvgCtK9+xA2ZxSF
Tbpz0DvDj4L+m8mMZCcq8Kgz1t1d0ICZ6YhQKLCRA9jeC1n0LKw8cVArBa1dHHYC
8JXSflaDkcwg5bo5nB6FZF1x5WrWgC2HEekOzE0zFfjpRnn5aLpEYFDcQAASL4Pu
hpu8mIXShnVU3RjJ42Wqk5+wrzCcW8oxZBehhZPHyDAAwEaLtACUTxBG2ygBVkpS
xaxZglGNrtaM5aERvnXm6m6w3Fos1Z/5Rwc7VrnIJ/G5+WmHyIN9uyAY4+A2UYi0
8kEPUD35ItpOCJ1JHDLGj/ItwkZjjLY9yh3lTpTsqPO0toNKnwNUi55nSAm4DWuw
2q3JRnqGX4Ipkq6qDWOqnDrWUnnY+7fg2hy0+h2DKHLqG8R0BNYO9YjxAvNVUZaB
3uVCRj630xq6e/ob4JFH16pq4PICttcY6HVH4XeNARfQDhpRIs/IIYrqatVtuK27
GloKkO4bhzJqt/CIq3EWms4tv+B7H5HEtYu5oMu/tem4wUXN7ix3PxBA2TY/VDO5
DChKKSgRSbc0hc2nN9es5jwWV+a2UyB+E1fFILoQtXsxajQPSS48ySa3vQkj4FCO
Sl3/0L1PANinZ37ZdPM2i0pLc1JOZ3y1nZR7IYpq+F41sqKC165pYYPLcKTSpsf1
YICdG9F3MPH5TGWIGQMHEVGrFol5xlVzqF5yNB9z1+axJn0SLmGz06V1fj1He0wT
+/QrezoPfwH6tQx+ToGz64uuvTTdJzQ724XUYAyWY2a/IWQak14IgRns8I19VLzP
L3wCKlFj9tL2Z3d45X6BXzfZW2Nw4uLIe/klPWNan3lPuMrBTdZQdJI+jObkJf+B
UrVHwjdWKZfdxxN+EzZUpU3aJkQgDEVNPPXEZTud7lC3/cpsyVKkdndpV5OR7cbv
iDo0rjFU8wxXReu/Rl09H43i0dfZK8LVkHlOgjZEaBv5ZqJGwahtoLTPf43BUIaM
cTelkbNMVpT3KHieVmllcI22sBA99Vepb8nokJvqv1kCRKFOI5CPb1VQYrCuEPPb
21JXQR239dCsHiVlS3BMjQYD/DTQweDE43R5Hn9wTrTm90hksnAE4Vr53av9i7Y9
97M3rQ7GmZWuunBZPooHAbMtb+MGiRyPVzII2mIomTnmOj5zRojQYP8fYdlvZ8gk
/M3lgKjzXDoE16pQ0b8mY/Ln7aRxweXqzpUjsvRyqR+Du99T7gH+eqkbf/ihcS1w
UetJY1ifOAzZRSuzsDdhMVpnHn4qSBD1OWiaw2UiZVuw32FFEkR+490cNc0DNd1n
1BsqAv+P33n/RIOk+MEKEIJnmDjYItIT2MwqyAEjrmDZWrJYStMDWVdXPcVMGyoj
Kj16BSo8scOkMKyGRv2nzoCM7nfon9SyPdeXT9Sy8MDCtIVnqSc41cG8n0xu3FPz
GSjLAMj8XSdF4jC2bbFN+8ECYTYYLNoyZ5aW1nlijzE01ShP701OwsdtHrU8XHmG
Sf7bkM1ZNcN22FITLUTlvtmZT2gpHhGk7DOQ9Mzq0OvyTrkUULZi8hwbdoh3Ez6I
t5vEvTPNeVgNOUazDoHZXIeeG2nQ05rwFCcpK7oLjufDLRXprFbt9kiSDPk8o94O
SRgn9ymRx4gy6mzrQ2HdRQAqXXbzFxQDVOWSQAzLO4VKLGCHNTFgNxOQhUkYRbzf
h9dsk9yZ+GSDoGMBtPEX6fr7bYplj8i3SfF5Oo5C2Y8XJ/v0eVxD0f1xwEmLSVDC
HBOKry2fuqkDqUfWShqsmb3nXbd8wWJun/cRSWzuapD8WuYyyNAxB9qxl3slwtoa
57gH0olsSuKpWYkSbP2dxck+AVfbs0iT3dpx87Zu78fgzqASloo3fPIfg4KAP+Tc
1L3+qYzgnn+FvTX2Cx8gHdM9BobdGUTxX1ifT0L6pLFWVMpIb8m33sJS/N9FJO6Y
7ES860vrGTZ8ORM3XlBiXVMtpkJGaxvg0Mwg3+YgQXK5VUE60DcUnWejPqriBOg9
F5giFzRn+0wcinRFRBxfdWDbidC0dKFr+xBSy0eEzoXvOo+hGBHIR2488gO2XKs0
pdmNHqUOpIQqJbFUl23GDOwNe3aEb+4WB9sdjClC/mHUikOEFitsYIoN4Jcq+coB
LxWqvJlZE2KvDEKpu30xBGkk0zqPTDtM4ks0nGcc8ha/D72Cst9Rs0oc/MD0QopQ
kB67tKfZC1+uYZN2ZihdizxQ86RxKRQTyJ0DYG65udM6uzzS+iMaAXamQiHlg2fs
cdgCd3X7aFXKe/Bu/3lWg+88attLpNPR80Xsfpf1rlm/SM6G1zVb6vTRP+yZSo1q
XQrwMgwExnZxxTq5GPEQqON+4OJoLsaRO6ccv3ZcsOy1Hj+At190OrBugImVqL16
DMFd7Q6tDZ8o8SonkWA5agNblk1SBwXTm/HR9T8MFZgcVIyDKP+lwk1/RC3X7vmI
Sv+ZAdg3A30/X7Vy+qg0Mh3riKf+wN7RmaOZgjW0XyGhc1FIdF/pBSacs29cziqP
fSz/riqSpQCd1GqMOYnPcpTHmytvwZHRPBSJkuD0J6I+nSiI2p71ypzptskorILU
sPwW8rbwpVgZJxauvVFn6ip2r6Jjl/SYUL/d/Yv1zp1NhKAz7hzQTWOqkfFz9Lr/
BDQKBUS9SDiMQlqT9Y/IDTGwXM58UVjgpdQI6YG5x//JacyOfdVrI1trYNtmvpzJ
Y1LZ4U60Ce/vHFUD/2UQL97AY8jurLLIOawQze5at4DWR5U9gnYoj/7ccSR8p4qt
8evzt6EIzuu7Zbczgtkpl+45TdWxdZY9vXICl002XDNps1+pUlqTUU99japtg5fu
wqVwp5wmWGB6yP2xx+PZTspfX10BimTsrklksCSTSH7t9yAG3BkKfuPvY8+n8QjN
xC42MJZHN0eIK2cReDRwd2I5tWVsMv80UaNyGtBK/1fPmEg/ohWqEEgRX8LDFiyT
ybmEekHbRKfRLNvtPSQ1wCtZhNXR5WpPfcwPwBv6Y740f22SBnynblWmkcKuVDuN
CDO1BeVxYDUjviORiCtYwqlAScb5ih/li0xeni/lsneGVmbAUKTcvYKxM50+d0x1
eicdDNVh5818bgAKm5ZSstnhgSwhH+ptWer+B096RmGK7LhRSK2Tk1eIfehnNoQm
+1lZRk5MAJ18mXsjSBLuOY3Bd1RLjIpq/XtiHGLy/ysxVTApSjHXMtxTo6vuxDcJ
0jKdGVCzp+DBVHJNOp2LGoTUsLYGE8SPoozUD4Kt8kMQ8kjFWycwAZps8IBY7SNj
0Tai82G4Om6om/qzM7dfU5kJ9JdG8Mzrzo0EwTyHiFzrIZfPpS2w8sas8UbNRn7p
r1/Xp6VMBwHoBZ28u75wruhdMmKDCB+vMmrl8eblGV/SNJQASi0PXc4A/i3O8Zal
5KKqcpuOsnkWhQe3tWtyj8Wfs+NwbrC6hATv0jAg3fI3TRl3aTxz5RlLNABptvhM
Vx/jYX6XD5XA+0Y5xGCqGakuZ/nA/hBbXbetuJCwktHAlsT+Sod4pEcBQWdwEf9/
74KkPshjJ3IErdfhOL64gzF8qdS1Adqh1VheqKXTVC43VlOTd832nzhxGpnEfcOx
KABYl11PWpaR1ZFBpETEzgiWvX0f4kByTv+6uB+hfooa3k96ELmQ9LIxUe+A0TYv
oYncq6sqkkRV28iWSRabTxMNXxgN5PGxxGGKAOX09udJDbIgs3JtaV1MEyLQ8zBl
Ab2vrMyGL0jNxOBlvZ/zYsLFZmIEhk6dCZI6r/pM08tonyvICHJXlpy68b73CrbZ
3TKIfpQyP/iaTCwcXcUfcjHRHWZrIrCG+mpeUtWiYp+C9+e8IsBMhxv0Z0Ef4AHP
dQ+OKHQYFEtTiNhtVP9LrQ5IW4XTU1O5allKUUoDTBcHaPsGuDGpqFHudOzXNJt6
5ok85MNEyLtisRUfDsyg+C//rLjqTSNMQWts6ogDB2maslKpav86mJ5xa2dALHYj
GZDlMjIJ0zXGKEAP7KNSVm9AXjrRFmIw7I2cdMnetbUAIs2zQcWUvTZ611l0a+Gc
c/CKi3FN42l7A+t5M/fvmnhhcOB7veFhUGrIOjxbgu1+b3+8g/ToBLDUr2hj0+Sw
R+6CMEvFlShZmpysoUFCdf8PUpfW81AGUCG8PQZLTIp4sHdUt/Pcgi8DjdH8NN3V
gjiHCs+qC/XB7uRVHMxaL88JV6I6h+Y5aqt0uPa+kMO71FqLGS/Q2tzg74lTELpN
Bmk464cn31QE54xnJ+Rrp4URsvClr4rCwLFGj9NFdepG9QSQ9vyFW9gATnieQhh9
Wbj/sqbc+OX9w7bdgyAr3AIEIV1Cd8t6zZhOSLNWk1UTimGbwAaKSTcd/snzuVU5
I/9q8ZkzYYu8R3sVI2PHyOgjXrh45V8K8zXKa4/mngN5K22I3hjcEOQlyqZUDZhP
ZgqoNdKByywGPrmSPngcGXqI/oJ/VSs9c2/iywx5bu4SxV5T6ccN2mIUE8wt5iFs
8qRae8WKP3vKPnrh3ggxRPyIUCVskW+kmO8W3K6LBVxbHYPyjlPWICMXLBhskrKH
Xi9mFL9JY2rK7JC2RBln+CZQSERLY9aosr/u5LZFV940DvruazqyhDaa2EaaROXP
RCw5jhBYIdaZSnrKsY9aflhTvFYtdpvXBMnWFGVW8IvQSLCXYDGpvJ43xebbBqFQ
zMBqSZs5donGoPDt9bgaz8a6fpJRndN8vmYcYPG0v3B43chj9ogZojkZomzYgmN4
QlPDJQemrpib3f34J8vTBtn4306FVPCQCqzQeRd9OyfWi2p4YD/NIDdbZnAHPyYr
jFZsq4GEUq0GpTBDRrA3zydljP0Ol3HJurz8KyPgypUF8GCBGHXA4RJUJiLM4LGl
PqyFxBIBLwoxlTfaxsJWwEmQ9O0Jc21fyStWlhOWEthnCxPvEx2UP8wnwrS9WbnZ
LXNIKA3UIp5wO9UuHqUldhBbFJOtho6VsIJKzu3X+S4eUgGvJTCeLOP02pik+L1p
GgIl3/oEh8VtnlRAd78rKb8sK6OsfhGVC/5+LxIhQkEXG11YXLs7vJ0aR0xxqvfF
HS0Ra4yMVXxURPfVlKSEQuDb7/e0CfsZIqLlRutC7ltU/fB40fFFdA3EgasKj5as
C+3s0frD5ZawrayWR1S02ALs/FPAivR18DH9fjr0d6BAGUF2tVLm55FdkliiH49+
ykAvYIJNiffiCD4h8sYCzH6iLRpI+ZM0/KbgN6KguAjOpCW5bsf31CJwmAXWaVUi
/1pIux1sqNpb0YBqoI5I3O8ht+M2MAVZBV4Tsy9lBBaVsGH30WKoVDmMAgWutXrD
dORS5PBK+bOksdgIIsduzUd4OWP8RVxP25OpFytpNEwEvwFvjBB2RfZY+hdSh1m2
Bcp5gtgfkUimRDxNh2KJrQgzxTUHCqYF9Qj2NuP8pr0PFwRuLmG9diEjOL4qnvTZ
BttT3+kjOmFQVW23VSM8h7WS42bS5rjH2QHoU19sGuXj4o+naGGZEPc8i8uxGkWa
60TMSZO76+5X4xLF6pvJzFxD59TIe3lRD6Mx9Yqbwk3e0VKzXg9mB5SKGBogtZMl
hLxJzr7ysdTcNt2kd4YGeRonmVtWLE4/9dXjsEm4tdmuUw/CxG+bBSS/OE5OUsse
XyzmhVFVnKp01xt4KCr9g4WdEaolWtUXdteFT5tXueQJmMHFzy26B5Nlr+HheSEh
4rUCUdJAlCWMnBNDtKmwdXhZ1exVMKWligun9XAYJlBn8mh5ct77oN4V5Uch1Hrk
jl3lzgLQZRGRCzrNI3BxKKjoooI4vEhxINllsm6uroRulT8g2kf3sxWRWpCogBAO
+spXm4aJyixkJUCP3tAa2ECfa1rpihm33YfrZSqyEULNj9JauHzjcGUe3rykd6sT
CIPm1h5+8GWmDlSWbI1M6HXKJmpNXrrQ3ATZxqLhGZrr3feVNS4giod6rxrSIJAi
MZCxWUX7+DUYKS0A97UsfJgVFF/XECC4Or567UnhxnIyYjlchGIo2+PIqW9j0ji9
8UgI5jxmTtrAPaDolbAli3piaVRf8H2rf+uudaz+zcoi0aN2fmClxU/Ggu3El6im
NkvNDkHM33AXJu1+v3Kv8MnUKTPK3t/l0YO5YD0uCSOlaH1vt42+yUpBCZPW9vW2
SHqG7lrketisY8Wrfu4+aRg+WCjF9ynFQLdSRClnRLu2mXiGy7krFhUE82VwJpbv
gK9d6yOILqD+Ev/eXVd2TOebmRaDanbhba7m6rJf85YoXtMjcd3SKuG981Hj9eQH
EPAn43+A/lOoDbzQqgBqyzFURhCESbjbSiQo/IoNVWT1d5TrlcqGlioFO2QuzSWj
nlwHUdims4ksyPQI+R+UJMgKLrIhPo2wtGeBuCv/Sc9eeYSKP2HQHbKn4PuWO4se
oIwtnFCNr8WD6EBK4Iru+G7uMOx08lpFZc7nIKlvy0yuUnwgcvVH8Ri35VBh/cNv
N1s1YGcLsAR8e3D/V80VbFaEwmRdmjApDd1zO0t6OuxKmrJH+NMCCThUNwK2DOFQ
HuRk3UeArIWkEbfMU6dyMiMRgVSxjfJwzTDc4OuYtAvvYafxN5JJqZPJAKyZnmH3
BkU0s8Js3pSK1WTGCcSkTWvlDAfSVUshshEMJiW5kx649Ke3LOW9e6oblYwJRdN9
TaB4pJ8/BmY607cmDSJwhpu4nmvaQECMui79OUQHLIHNX7SbPWsiiD83nxZkrkyp
ZQcjPPh1gT65UgCXeiIpWXpiFZO9xCR59qAXcD1RmI20Uv2UOYHXZTDKiEB1rZ/N
G5mlIPus8UAy97OGQp/lll+LxO1jWOncJz03N4tqTooFB8aFWS+OcWIGGQg6lt+c
okrns514PyDCQEFwc7unowU063DLUWo+I0QzVR5CfRf99LEPml1ogiSCl1GCassB
afNHfNbNV7Q3c4kwa1463qK76vF20nWZjs3uFevVDIYSu5csFVe1eSC88sAhCf76
uDXLG2PFDExuF5sfDXkJ6ZQx5m3WArMTfdJ25mU0RmITF6/pP7Sy4LpCivikdLKx
kv1l6k/ZHdwSTkBfT4j4qVkBneF/8sWAtUPEUV0nNFLeWzLz1bcXXbmJIQF0/fno
WLrcD5VxgWMfAYoBfx4RfJ5zvAyTzb4rg4eymSnzMEeTWtncsaCluNJuKDX+EROS
Ny6UxCE3wygGu1Hxgm9Bs1PiheUX8Sm8p+SfcBKDcBe3bFwE3lUjUOh0ay4JqyJC
+Zskgm14W98Wlxfol4a7a77rJzsPvUziHfwQgPdoSLxqnYJp17nrSdORbl9prK2q
XgzOmpoDXFm5nRUtSnNS/4BfOSlL5j+qkR6Do1KXbqMaRK+2KgM1UvVZMVpTWe7P
5XwLRof91FyrYI689HmE9ZZSPecmZBDXsw4OfoCKPBZcCS0cnF/FQYcARhSVe1K+
ixPQsCC8+mSA6g9mopkZLX8w73/Z3kzNvp0brwzMh3loQLbBn5Dl4jJy6xJvisI7
b7gKKNHKf5tszkjicgPsEZF41JaFOi0CeavNOStiJGXUjmydze079BHHPmQk8viD
3a2FKUxhvYJiN1PvOaqZn/ik7Pko/OguR4hS+r61ew5AI2h/PVRgY+FC9xHC/6JS
DE8zDOIiE/S4GlhMvXlNjC7MTn0qznv3yn63GATk7x05wTxtI88TAqIBZwHbiSXM
cRcQfG5Wy+uKzplkXZuRsDPKC72hQa34QNih+8OUTW1EiZgFDWNH2xxrxsy7rzsu
JGLNacdWPoW6Y9zK8/2UzCCYF3K6rImg31Ey1TN4uBLgLxGB1W31EOL8JehQAUai
bodlDiOh/5o/ErB3VVncpMT1nB9VrMhhILHWhJnGRdDSrJ2r61q/JxRZLsRL95JK
P0LWnoOSsrrUOAG4Z3aVs31ShIRGSEwvX9VqExYL6tdfkZdgQpGtKhvGaavb1teY
GGmZtbHUJRv3yoGRNdMXAQf4SnFTtc0bB8Y7pjqKTJUGzX55a/KzYzQk7AQiEzNz
Qc6JP9kg+wNFWbSQu6w/srd4fR7utMeXRrZeClivFy4bfQQHM2Iq+eI/ElD7MXNC
81PUX8dPrsHKic8vH8yyFJBhAbHxRuBhlIQYIpFqCoPQvT5FWd1E4ve3gMgfYJRi
2rADrUzlQ0JVzcpMmaawwH5Xz+TOhF7/cFlCk84GbGs+rBQQ8dWylXCrbhcXyN2h
IGxcNlZXurDOgWu6pxwiw44VZ7GtyjBMO5L7rqIDogo0LMHskxD93C++dfyAGsRz
1CoGlSpNr7er4d3+tEC07ADwpo5JmLhg5UbWB0QVoNDqIGOdI0sdFYYL6zbUWrSq
/OH5vqSh5EVzCJgUgEpVtSkyk3TUC3cvzSNamD88FhcJ5DCBV9FYFOAsjo3SvJ9H
gEnx6nvTOPC67i/A247ZTlwjDnfsWwdMRIv6zUPuYpuiKj3XfNU/JuFrYnlU+BAa
Y0btxif/TDnQt79Ts7skETQF+Z12oVeEbSrxceZNOBcPBmwLhZio8S/Hx6MLOJEl
vijd4haKqezrCiBbMATUUA1gFOkgutJcxU8vgeW97ngK5KSueTJpxJ1M1hXpBuMc
XrPgPEvEqf3+UgxK1P9VnEsvq+Rpuudge5sSWG1kJww8BQsdhP1k3ogwcLeGEWmo
T1BLi3L3ToEQ7aMR1RHzj/J9ErSP8Nu3DcGyz7KCuwD/HOR8k4bv3RiHX1GDNAxC
YBKZNxiJ93M0EXU9my6/zobbm2ZcA60/ct6JNbEF1LItLtKubbUa/qRoukbHT/6m
xTDvFjBWlOiX0SGtW4n7AZbg1rMcgVT9iHO8aVAzXGJ+Va7Wg1juws5EYkBoEXEK
D/svpWNbBSKg9SiJv/00qGbM9i/LxSXqfHsLwiXR0K4r7cWCJT1cWdvkq9glGTqU
AI8BrKPb4ivOyCMNlO8VedQ4jQlMMMUCRMCIj/T4UqvHKIMfgCE+H7OVUnk9btXq
T3KVeCPgTl6qDJNMh1nUXNlV6farnHcrKoxLoKza03IlBzrFKl+WsnWBunky9nVO
JuaK8AO/AIbTuK6abpC2NVbxXYKzO440YL/p982axJl3fmX8wG5XH/8QTqSyenLm
BvpcXNhQqRaNiOT03V+qdrtyYSJpPwkYhjOjbY/V1hTt4rKzKTcLDGipGHYSb0UX
DBhiDLiJ1O+Cw2AFJpfP3Xe2HQAveRix5UxUFWvO/sSiuDThKGvbVSGoc5OWkig8
jlXwg26fFU2XXcyMon2XvXt2QKaGkCd/COKhNUSjca5zmCBsiq2k8vO8+4xXzhnn
9LD0ADQOHvmcoWbVKzYE54ZsO2B3zz/sNS1gsYTXwNwO2X16EflWTofdjccXM4RW
qB2JUxVBfeH7o6638OpQbmJAnEZqQQ/Xel0pPBd48jIK0OZKwhndvfJ8ExZ7Tk0s
TgqkK6XGiMHl+Qs08mgoYpLgss48+NR9TKOYe4zOALV+Dj1Q9YZDdtG+aqtbMD5i
dXqY0NYI+JpeDlxYMF1NtvTvu7hzIvsqgGZAUvCnGgZNB39y4q2Bb9/T7yNtYqTR
7SC9EB4keEVjKF4UNI2xicq7eU4lF07VcfhMDx9vm05wWEKAeYQKjspPWMERNNdg
PxN+n2eMsxmnIvV/bTs0R9usbQi7GuMkc3p4P2RNn5d6eA96qXezsOOva4nyW4tY
cDj5AWJi3DF2L0V6lcoyMLy4C6Ua1YE/J91/a3+bP6YkdH8UEjs8wOsLGnToHumt
no5oOITtbxq7+1kZ1QF5EAxDMQz2rbQ3cIJ6/yo/P59LH09FHcOqZnEbPdjgtwpx
3n13hTsUk21cU60IMQ7KpOXcL9uM6A/FTGiVWL7NAk/+TXk9dqGZkg663W1Hziu5
ypis5be5SYyC0Os6oaTuoCrxHTWzNB2nNdIIPIIduyN6qimqtthQDpFSXiG8Vdr0
0MRLFmEa8YHAgZ2jkUnGd8gQ/nQ3XcCA8+tx2pb4P00Qo5PzxJhj4qoMAAFu3CGU
Dz3Is4A7Y3Xz0SzBMMz22r3XjP0Gkpd7sL9IgLDFjsLoDhqBF5ywA9sO5JsEHyNe
g4CGyysS6asxPhAzUj5cu9/ZYw7NRPclicv8KHGcWeYUrvIfhoWGfutCGyPvkrSo
dIFdkVJV7LguGYzf4hY72GJUT7iAadQJ6XLYER4rDZuQtClUkC54spWZO5/zKOWA
oMZbdxf4YollxOv7/owMTS0U1jMg2FvudHZ6sI5EiGGwlF6a9D9nP2bwd6ru5kPU
YOjbLmjvSFusC8OP4h7js3Ji8IuDSEIqRYXwaHnwZ25HAwOpUxAbwNxC79fkCQ1F
z0q7lgJXFb0/QX3WgP4gzw0ndnaDmj5ZkE6BgawWccTTyl4xPyvcTq3BzcF9dO+C
FRjS1X1XuLbR4/xtn+Q4RpjFCfEXzK9oRs6oV5tpANkRrSqIjJiubF3KwKlJUKyg
j/RjOn+Rl7hjhUIAoJvmg6+gCkm9QVPwm5m7oPnY7ZYwequjHH8CLB2Pa4Rm+Wch
o3IbI4gzhm0vgcHY3vETaz9Vpj8IQJVYFQUHhsXAblfN5MWyUjE8PhVqBGfsO39y
QR+IGh6HRxu6505QwL7r5RRInRyvAUv7HMVupeljbED5G44Ag59/63ATvn+XMckm
L/jPNWzsRY2YiwsVDuFVhislk2xowQmTgsQ2PNynNLut0Wx4tuZCwKUQMZHYvr4X
ULFPtBJHyFkpl1uai1RQC5PmuGUrT1H58xRpWpFE0OjKlPwEEy02xRsehdQgTCWb
0UlRK4bIMsEMqxAcf926/xtHhQ+1Lvvj6ufSAy1l6324J9KJwH8sKTBTKpj1HXnr
ihGDxpHGGWPpqtClkU/E9PsjLb1bGiFO7fQLEeNhA2+5A0WvNukolFvxaz/PZMeT
8YHWwiPQUAnrl9gD28ODQx2iVeT+2s9S4mHrHHql2gQcO5oQU7ICzttA02TVPFwn
cy/DltJ6b9YC9SEDLsMRgLFDTkAgMi+kJOx/PATDFxzecWht/D5EuXfkwBvwoJ5D
UfK+v3Twwqg5dhsBZyBPE+EXmQG06TyfgQRKVqrMckjyN+aNLjJbWxBRpfdgK+Po
42vT3Cs+Ovz9abI9gk31PuBWHi/S1AQ06RU8QGFTc+kMKEsVJzNwygu2qeFgm/LC
e1r+sWtLorL2M3lU0tEy7//GN8pO1aUTNX1TKtRf7GW0M1nsIbm/mHETvgH/Bps8
bdZmnnXQvdjXwQTTsXFUcr9lsD3RLtw5MlpA351igpUMwMbU05YsbsV0jy4GUXwT
xKHTDiL/2KT+W9AtclEJ2raj+3RYz6eYsk1tPxOXBXf7RhdMZtk2hnBgCAt9lL2m
TF+4AD4KtDMpk5nG5GKwKz+CJcSjfYr3M74yk79fsGHvPPDRzRgDBSvlgiJ9DYKt
51GAbNiKCjojNpC1DoHRcg0y/JLInRaN1++Y+yMcSYGXX6EwWE/oA2BKDJ3+ckeT
5S9Wg8tjFCNvYcuubRFBc7cO/h6k1gv9B4F997g26jONrFO+QiKFgeQ3E3aqfN1A
RGflyHR0xGiXHG+PJRURJJkk2wJ/r69xXr1nbH+j57SWwOGWjdzhMi+CqW3MgQcX
2zBYvwAAbfVMig6tDv6FVtO+SOetNZ++7bDOBgJCVgkFwzWlyGVd5MFCiqM12TjH
cIqPYgTalGT24xcEdtnr2RR7qbaBQJuDMTCyQvdUF2BcLL1lrwKxjpfbRNwOquE9
5mQGdO8+JER1s2WiWg/Vb5eMVRGis2B2sqL2eH9FgCaBGRa3Ue3+4o9DS7DBWW8Z
sX8j2Gk4FaxQvj99voxhaN8ZUHq8/kjQxWj5EyKcl/rwn0OYO5GoY3tEp7ogtcES
NDHfRIY4iwecUhfUkF2B9pkWqDA377L8BGjKtXFS/nHkEU9cOe82o1vf4ssfkO6e
/kpd+OCYXqyUg1NLVuMpba3CyFG9OgFtQc3rO0Ha61KNaapY+iONV3IfGlGPErcX
yW3WuZ+o63rtoNSnPVYX/y9vxGujlr11Gp/aEffLn8QpaJtzWNIspjQijjRw9Agj
z0TFBksJQFzOaJhjsxHUy4ztRd/WKytNo9SOM7M4gglqxPoWdSAaGj1Gg3eK3/51
V2Gefb9wvF0eLv6evEzjPQQXbGUJfDJwTCO9O+R+YS1Y40f6JA4FzfYE8wjKvwPq
CVZv3BfBKlE6SoMworBoctM2wtBDZRPFJ1DCWmrqN2cH0I3fJIReWUEcOsQEq7X5
h5KDxMPJg+h8F/q+4/AK8IEElUD3sZ1Zph1yJZx9ibMVwbXjQHe78qip5mqLDYi/
LQdTOCUN/gcITthmjM5jgyclb6LDmn67gc6bFjif4PAfvuahUjPTUCBS9keYGD+p
mW64CjDcRkn79UeD9qePspVFyUvjubzG//wUTu1oCEX5pVPwOYWQzz2zBx6ZuW9b
8oOvNFBgJUjso0cz6ofUyk6O+5XaG9m+teu+/3Qmw74btLnXKzowmHvT6SFs303v
JkMMhAHeRTBdR3CktPPTrMsO9QbF54aKTrYtVrQIwdca94F2DYTctsOPgilEGZDc
Xa9rB9JhVplQsP5PMZTaB8MhNq4qvk6Y8/I+qhIArOzeeHvEp0WUZiL0mDcHIU6W
S8DS88fSMQGkXdOJlf2GiWL1aTerJ0+jAYJW6hsnTsPTS6Vv10DtKN9YEF4EwZSx
RRUj1B+ya2/lfCHpEAjCqXrGno1x4LB97xcbf23ZMRXWgRW/0AXxtH1OWG4yldak
LA6x4gCc17tQ6aE+/FYOOFduP0KKYylNvxe2Ra6XMEzP7mLcwTQyEWEa8f/Yjtte
MGR/FLeSmeFpLwAVQQEO0TWjFxNXqPbA++6xRGUgAvPEsN/Y4/PkJHRVbe2GM10t
F/YK+Vv2mU/OWvLPwMR4ZWLeCUxbClz73BH00CuJxU4W2Bl61+mc0lMyNnF19OUE
CJzu8cbn6ck/dgL29bMat7kp2vpmikRWyRYW63Jj36XTczvY0TMZ6aRA2nSOSOKq
qJzLIBQK0AEAh1KDB18G1RV15SBq3EyC8hQNkxh1bRld4YwdAAFLT7C8B3ipfYzr
cIUtVCmXm7jTImmOt991/qmBKVHhq23ZmxzGY9YkJ6r6QnEXC1P5P3hiNV2eU6Hq
BybisN3LaTiVZvTVHOZrBRnWqD4ocktlRwNGS7fXB1WBVhXPCnvlJ6GX0M0iBwIx
PfbMl+q1gUVGxzQ3DQAHs50gRzTIURtKJZFYJCuVqA7eejMYzwnGINzGHHisRrHj
LQjNA8/eeCfuX+EvMFBDvkBPQADwUpfS5XaDD7MbbxKedRzGU2ASPtctecz56CGo
m4RaixN1BrAD7bco4NKt3NFa+TAIgxgVqswyyQKsRCwg5xFjfzu5nHlFZLaq4UkE
nVt863sJKk6cw5wf2/RBMm2XQorv3f9KU4XpggOFnEPvQI+hSjnGQ8IrLtNaxepT
S75zXYYE8OkrieyS3eAI4gJzXis4+WP0dAE90L5Ty/XTaFDDm/iCCTsmSfzX6Ypy
Co7mow+tw1Orf7YleOWcKVZxQzaEF7aNax1IpEsFhwvtREKY0rFX8IWaJV6z5/g8
8xsRS1Wb2tE2RXro0/0ngR4Rtu1M4nXbImzqCam65kHZAYub6O4LkxrPWtRoKcMw
gyju2FYemf31ixIYoWJ7uMTUzQeu8iwjIyticnk0XdGsW8ye11DF49drGJDvnViv
qHv82ZcUXkiH5V8vVI4I60JVeY1p4DKSW7hK+RhR08O291iAS/7RS5jlvvlTotW8
oDi8BcR+Bwzh2mDkixKx1r99qYRtwUaXgRbWQDA5SX584VKEF73aY9uyp2kcQtMZ
QubbZJ2NvuLXNzPacWydLD5zEzhKAt9JnPu21n/YtfIsSs0JSf8TqzbTzm+qwFKc
n6BlBaTeqjRBun2hxohT+BHAZLJdOZg6EgZxy+ijeS4vVEroGV/wQxt0Qwh4QLp5
+fHU719bIrZlbdbZH5BcpubvSnF9ynvRlwfW2w680CZFQP/U5Psr14jFhoie1hGh
fmWGNXfLPSEfy/j2kuP2sDrowjvBxTLubElUthFJSsOVg1oL24BXLK9i+rwjbD6N
JOO+Ea4BAb5ygT5FsMSLES4shWZgolg3YSdXASOXbaRcQ+JkSn0jPQjrrcfZgU8Z
x4vFcNNdfjlbDVXuHHWw5g0j2hEeL2OidsE3rMcpuA2DkFESJuZA+cB1IHI2/+4v
p5mlvEHu2mShAUZ2BX/cZuXQufq/LPj3QKkQPbtwUbxwD2jmz47NTI4psCL7grRM
KVMLssmmDRNeStOPdcIekvJUkw4UmDG4Smub/2hJWu90JEbmMTc1mC/gLh0Ma/6r
e8hwhk0u2e5ID0GNbQj02Q3iDKemK3GD1VzWdl5srC3hZ0iHaSnhgHmC9UK5fUPL
gxToUg7LvN4NqC4EkwWLSpgMUG4WGCYchQQfmghNtoza4CIcrlQyfN9QzYLIUkIl
VZ3cuK/65vPpaU5sBn6D1CbER9W1MxYXl44NioF1vcf6f7ySKPisLUT/x2fSp7h3
kw/SXJbiJ9BKu7Yk9bH0dzO51kjVpRbIQpeTCpcB7LeXNP62Mv32sbh2BybtgHqu
HSzjxbaG8eLlyNcgGaXtkeQN9J1ZW60J9NsX2UDQAFF8jXC6XD3gFIWPiuk2L7dl
qd+Z7qYuDGlH86bkpL+WTDiflywaU7PKz+59tkXNR/bazC8TnjhuOPui9w+iI0aU
eUiyrdP9rxgFg/BDaRI39NyvNG7XP3RGdNph48DD+Cm48DYpNM3ZFnCJldWjRnL8
RqWt+ZtztClxjmtqQwzQY3cqBjiGMzdM1ZgbKmbg8YIsW1j4qxkHN66LBzWAYnXG
0CB6WM6965pOBQfuGQxM4+MVfLpv3uEIIcHMZSt3UnfxFBQSacitET2UU6h0uCZf
a3QtASD9eKvtgjlLzn8LGFXkWbTnysBYG3I+ZcrE9RliDPWAd93QVkXZ5AqyQuI7
iFk1OZ7gMnwYCycSzsYkY/GMSWAyoEKVJpufdVUKb8b1hGj0VWrnehnf+6zFvcQL
1Q1Z2i2wO4ljjrc/TjBkdsVkgZ6YJ07l7Ln7ic+wnL1iiKPLigII1MGSpMJNIbYj
uCqL2axUBt+wFkB6Rxm7YCbFSCducZ+OsDC31JlPRglDaVLRNzpwLiJukAgIZj2Z
vj5GWTTjur80uZGYjwN2dz2Y8/VA5RBSylbi4jwC9IhmMRNranx28owbMj8O++3l
x2Ui8wZnBXH8O6ntnL/x4HG9xJEzh+kO0yqz5dCCeywmlUht9nmKACR1WEBJbSmd
LKWvy21V9df0djaNQSHCaPzr8ZpHVgJsHroGHw2zMwu+8ErMYu/AUID+34Oycu5z
JouAvfTfCtdXhPefmbm6fmHM9HVZwO8Y5tyhOvHeSmCiCk2ditjmjpRM5WJBcmRR
fHcHe2t9gs9w/eUHVB5uuivHmAqa/ilI1no7fLqXX1IrAzDoIpNGCycjYK/XziEg
O+9FuucZgF1tt2/Diy2VAD4je8TWkDOgB9+8JuRBfGwDX3lRFiHn77VC6je7tM/R
Vnaeq2i8UMTce78ySLaRZ0OprlnDHnRRPs9YGe8boICF1PpRwP0raMJ0jhqttCkZ
qXZp7RvfglFv0N0qf7mZOv26Ljw0I0B3vpEfnPhy2PxtT55olHjm+WNEm5AlMoUp
Wu7TWfcZYwaaGjQaCHU11wubACwF4rVVsRHMH1eidI6oXsHNaJlh4DEVL/H8K+Ss
/DTziix0RUwNAUyAz/LvbtSIlQ0pe5CyYP4/aQY6LOBgijeeLc3hWztjVJGs7dcy
6QCvatDv94mANVIVja08nZVDrvDCOiddCqUHQiVz7h/vJFqGfO3FiLqxss7NhOw1
3pGe1cKgvYoMCCGmxCGkZTY4gOYorNyJqWp1Tg3YyT7uwsKi3dyj3IHQNDaz2Td7
cgc0n98esQHV1oQocieQzFyS763VpHSRXcDbW3S2aNRwqH2imeEO6slV70UHUvPj
x/lOkQpv2aKkvICwQqSsm1bRFHaUew/mPgMyGl/ftr0QLZPOCM38ttMMy4vNx0Ts
OzLPYNFLiJR2yEIL+wRSnZisN0FOWLmbGjmN9XlKhXoxq+Zqa1d/61QXn9+QQTZd
SH9rWF+HxrMe/o78R/tYHaUuqFiWJ1fKSGQYMAgDRiise756kwk4cTEt4yXMsT8j
b5DSSon2NXNCrdfKdi1t/puNmZ7hhfMnJURwTXN+s+y/nLt/txKm0J92nTXfurHp
EAnBbmCvaRRBLmLsdw20H8wKj7yRYnCr33EhWQ9QVta9JcWCXDjuD9OpUXykno8+
iJSG6qPsevG6b+YQzrkl4/JhSXVsDHNh/Fct2oQ558Qutra3gNkcL8dZNvmj+CYx
yYI/qq4BnEGa4fRbRc1fOxRmjriC0XEncNaEEdWnz/5aI7Hwg2iSlCjiqc/2zBUy
tyrJdst/2eB9AIKsJp1HxLqKq6dalRgtUQJDjY3R+9KeE0pC8hzQz3uA84OIfhkr
Awebcn6GPbELtmKLz486327Jud9WvQLDm+z1e0cMtQK/nQ04Gaald4FeXqKUT2W4
WygFKdfsXmJvCs7SEj5nx8D++g6PsYqvSx6nAdMEzXy1/DtYkzW9MTptQwq758Uz
bBdK5F7jVBJ5yqz65q9/GItVEFEyKdzEcAtNVk2t3Bei4pwmEQlMXct76cPwVf64
I7xF/34hFItC7pE6G+OmKiVmidps8XfuQnE9LNC0oCOleRrCJduDO+DclmHDEJlS
+JswO9A2sQ8d8yMgVBxHyz23F1mQhUYV0qVqK18MiGGqKrZMt/Ir1XhFJnNbseMH
lsd/2atQexm1TocZdyd8hLKnvvvviLeC9GXQPEp8DXxOCYtslgp4GtBET/IJ1/RS
NpA8WjxKvgnHSsv3hr0o+JttqLgQyatoYmRgYgfxMqxBLIrRwxLUTH5SNC4eb5Hd
o5IcGdlReQkAVbB+31uPmmvDDxLzKS0Kab2wgE0X8XvPwp1hw5XAKRwdK17gElf0
G1xVDq9bNpAcBjpMVLdK5f9u2OnYHC9f8Zm+X5K26GLDP8z6fRaiomrCL5MhfBol
FTOMCiRNEY6oHixDXsP3k7mfTlmHj73NWrimCVD8BOOU0c0bOA5pvrq3EXIZYQGr
ond31JsY6+rlgxtMLcv90FH+lkSUwI8EGZ90LuGUeAYCeRwf4xgS/uIJhylKE1B9
O9v/3dDg49hUSFTE7D/cSVD3KnNGY8+iD1KIFvPCL7D70aNlsp/XlAHW6uJN7KHP
Aei5VrifpL66riRKrGepjvLUTS3fa0siKCsC5t3A/evcZf53r+84n8efloYC06UJ
jCMszEiLSixhdFIW6m9jLw2nBlKBHB7a/9ox4FFrDWQeqz122sbvW6VUZpwWmPct
syNAGWJgwrhsstKER6e4/U9sbKxY+g3JwNRc8Xv+v3JMcvDkUqbjyZn2QWEsdtr0
6I2BQf15gTmeRyx2ZTIPnthxnhGsYfZMZJjBWrCwJJVC/NKzrCwovOmsFwl0fVvN
pi3TmPKGhkJgFYrNcd51c1MW31Ko/AxmzzNjs/bkJdm7yckTD6fcZyg//yN4wmNE
ONd9vetJi/35YwVQqUk/XajuhbdShB7imhLZVzo9tONGEzc1cHrjV4bLXZ3VM1SL
crd2+p/588VfcsTGCh0pCsnj5eddp/mTjOAUJcQNGeSYxftS/YbNDPHS6Q5ItA1d
Q+yVLMeLd2Nljp4JVMrWXurswZi/gIbqeZg4pniqFsx7P8Fxxgm8uZqs1OoG6vYR
ysN6kccAjfoM1AsyGb/sdpyECoLSMvtF51OOZL95dEUHAGVwiH563GFUJ722G+Dj
LjrCTooDlwO/tgtJikt88NttDLjS7DvpvwMVljzWAo4s6uA407qgNltVjGQtciVP
+4jnV1EMp2CQbzxLRekCRg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JGjNwMyhfwRnd/5X1gEvR2jWE/WgKDLPUIQJ5wJsijtIiDGUCRQnBPko60JQO0p5
aRrPSgsXsSjlEBrOsca6I0533yDFsZoMHreIZk2l5XqjCh3rBEZFsZvZnc77ZG0z
mAoNyutCid+dCQmT1Hsc9nMT0BH9UQXrpDq6J0FK+/WMa/BjDu17RZHTNUhYcIMq
osR+78FPQL+ToT4cYrJcG+tTcjic69sUw7BNIb9hrpLm0EiVBDNhz53vzUv0ob76
17hVHTh6P+Az/mah0Wrkw/C3qCqJoiLGEQr0iBQur+kkoMUgjXybGFScWNMXUiYr
wrVDrKE6vN+UPTPg3xxvOg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 24720 )
`pragma protect data_block
n1LMF9Dyz2bzmDjur3oNsBeZqQmxmYHBX/x7TLKltdP36vhM9j/ANmaBpxFX3JHZ
YpXg3f85TRSnKMvLPW/OWzdso3Tsxs87L+CSEy5tAQ9JBZUDxw+HwVuWrwdy07YE
oZF6lxI/5pIPEtkaGVAllEDdUdQEpUmDHVGPI2vQeiyprLTrevhSA9lgGYNJQ1/W
a74WB4USaNTL+jKcnJkSU+tvuN3MGK3DDjndRzsN5bDAKv8WEYMTyHkxntuXd3CY
ib1H+vIdtk8TMkWGKcDIPnQfiE0SueU4gEe0PS74mI10VBDmyaIJf1vAEJQ1s/w6
6L1xVTXC8O0nG0kYTckMIuH20ZHv/W7fIp6gTJtYfGnO8eZ/I9KK6al7YTyH+JIn
vbTujknu8IjGXMHLhefR6NnqZdn+KbADvPdUa/0ybD03rTSyHajIPI52YucziB4X
57LqRdC1H/Jv4z0jBvcfuFjEG3NVUGcX+azljoX60SsSu+ueNrTe34Boix33sc/Q
xhrESjNnNczFCHSCRe47TReZvBV46FvhezDJbPBXLKe2XXMKKZnKhDWKXmRMlhbF
Bw1aVaJRuahS+2sgZftuAkAOnBWh4o8obhcGlF9w5BhCz8pmFcIMHFnFrfGuMHp0
MAmILU0wzt23IquTibB5t5arH+rXSn7Gk5Au7xnii7S7TrMg0rERRkKsB618AXwN
ZUPJOoxb2vQcbauufnK5hvP9VtBlNpzvgd5YxPD/W6pp2fTyKQWjWq+iQrsdH13L
0gp5sDDqB36wl1YUisuZRthH0UamciFkO12J863XXq6AKXl99GKp2V9elSJ/dEY6
rmel92zY33rTXGdtx3xlh3vT6N2vJZw0PryFPtZ1n1vqyCEZgU7AR5wbcPuQwJCE
J28/27VmcEZ7zHrVH5TTuSqc2HKUEc/kRVWsR1H7F6WQo3hwweyFnzwU8V9RjsLE
u9R/HYSXQjdA3po1DGxEbjvlt+sp1JBr09+tpIypZWGqp/oBNl0yoaYaYnQSGQLB
uNU2ef+2r4C8G8zJDHerVrB6O/gk4h6/vR7+rhInBdwtnaY8KntmBX5DJEZ45+D1
AuhMY14u75nVlS8W899+DQvL+1hxi3BJn1AHC+XfFmMOUG2vqMvOZeuO750jOZXT
Ms60Q0OYrFExy6KIg5MLJu1UDwHL+yeKQ+eDGRl87OnObd1fd+GBNnqFcI3JkHdD
4b/slZ3fJo65T5sp1qsG0pI3yKxvOAkHGOzHix8CInUcRWPfO4I+Fplm7KHmx4JT
fRnYdv7EGt20Vmbwb8mui4TuISJYlI3ciNKzh8YAbS0UR63KGksxuWcWGxOoFxXk
CBi3McZcGZIGg0EPMNqa6n24xErIJgxG0M8H2jQFaGRWJcDDtX3Xn8AJnu3gtKgf
RBX0AT8HQ7hzUCSaOVzGfv96Si1PjQaaOk1OGZpWyQLiQ0EA0fT9Mq4zDe44nrXc
J4HZtUSv96unG07Qev/LVB9ga3DOLranBJdAC0y6F0A2JqnFTaOObHkgyQzM2ETM
RIeQ/URONzC8CXH4dEbnGUfgxaVKAFDvwZZD6qdMX+ToToAQnoM88PPr6mxVYBOn
Qd9O2fvv37cAViTVcE7F4B7XQl85dE+Fn2Vmdj913Haeen3qgzrwESWz/grehTWo
iw90ldh2k2RI/bHhFqDbr0+cjyvWf1cAXHuO5K8qZ6gXJMAI6o3h3J7+loE36jN1
vrvXgm7oBERIlbrOMc8DJaXUryU6IWeLCzFLS1jnrUI0l9RaUb38xlrWiKeo3jgd
atUdiG6cajdYgZrJVvVKALeM7D5VaJ9piTdcOHFyfd9o4NnpX2O7kE9AGFHlrxke
fgZRm/8Tnm+O/QwkV/DiReOywpoH4x++YfwRUghP4I4AKB5juwCPxCTsnU2FhYyn
mEwGfEmVUQTtREe4PD3y0Agip+yckmDtlS6DPBnwaijiKIE01IIlCxGiB6uvb1rV
8/zRYPaGA1lfGWA63rEjBla5KMcat+ogptfWhYOAu8erzGHotWjHq1VJMmbtKJ//
L4NT7epFVvDDAMtaSWrizvR5HDi7baCGYs+1qNkU/uVYR33K0MTEyZ4faTaIyWiH
ydhlz1By2xXZR7z2e+f0xYTKqyqWK2lIj+jnthbXPFWAg69mcaZRX4Pj6s5/vA7L
80lYG/bYxrfsj5IiKp58zot3MvS2aI5YRdZuFYoCW0OVGbizdyePHgj0Rd6e+Nk8
71DR/vM3/yGUxEsoCSnaup5v13H3Ns5ejIazoo8tkvK18OTuSHS6jt3JmWouQAqs
N8sIPrRGUMHTTDgPhwvOLO1eKNdNIZcYRf8veJKds0D2aQTLyRNw1+a8MaK8W3pu
1J5hF0QVx0GqmxAACl7DYpd7V3igRLjfeukVVfNS2ZGqfrUVguD2oQLiE2eBGfXf
VYQ0hGXpD+1L/5xtq42diN02EeG1nCnpgH+PnQ2XT010R82R8/ihdOOLip8IKzsV
odVtYdAM/bCI9fk4/GU+FniE1tfJfHeD2Q02WfmlMvxBhwx588ahfRIDRS22uVsQ
9IZUNsqabE0fhh2cwC7IHNeTcIbMGVBTCvOrHrR7LyRQmdH/R/brYAAXCejukO7A
4MIKzkdOTsNOisNmh5/zjUoTc9rg3jWHWBDosp9PrsEN1LTjdRRmuSUmh5aNNjXb
nZ55IMME1p0SCnomLCgvpVaaJiOXopadJ1VF+g5eaN1xcIEnB6633iPZUojtwm3l
sTbAyyAhzpa7Ko8ZmMqJxo82fuapyp5JonBD66LT7od59ecu8f1aP6uc7I1FXMZK
HjF3xSMxQ483VqGxuFN5AcykH7d72tKRZvgyywjDxsCXAomPqEjB3vDk2cyXdgBy
oghitT7EoxH+eJJ8w3IIcZ+Qim4Boy3DBT9/Co9lnqioFpjkpALbsVVv1zgeU8bd
VsuVjWBLL5GbU0gKah3KOy/BQa4KzVlAhNx5APQLe+Ws/quRtDUqTorJuZvTm25z
HXT/6xYbv8sLJjBVjTxf/YqB2iX29YUGXP9PY2YHRgvv1mMIYboOizmSivFGdlXQ
PVVPGuSjhyAZZVxTB22awpA7qL/Zyt1f60o6Knt/fyXwmxe+k526Ob+fvxX529ur
3HKsyploY0a5OyJVF/5n33je9Z/49b1gyT6U80+m9ja8c0IcXCSRB2eDjrcSh20q
vlR+w+iKuV8dfxWQbIfz1PFgSVJ6QpKWgOiwFJq/mKeXVBWOWuoeCmQ7xx71TB/7
4PghYcWdx7zhPPInGI8CFVJIsC752TqjehR7vY5Q7XhQI9hE4iahDVRpy7ROo+d2
ATZDvXCgc7FnfbH5WK9Gibcd914xvfg+t3IGlYQPyvYqb2isGWgLNmi6RlndGWYq
IF/ckwAKO4MpuUmUqH5dBT6xkIS6MMqdNvIQ3eycpFyxmrj9NiJFd/JSthGO+bx+
k+SUCkdNC11w0cJJyw1FY2Jo9ihZvL79OWvQusR2wUhDd3BmrYcK5+qZ7P27D6cY
xbns1ELdy5IgsavmdgUNH5Wc+gnL7HfuYx9/6jlSK3NB41PB6VdnvJmyaaxx/f+Q
ouPVEQBUEdKe0lVdt4tpeLS0cbfTaM9Y/Q1molxsMtZfR6wv80J68JMfGyIQcN35
6t24eMTNHgleVnIHFoHeY9kkPgXVeMztNTjj0as+AFw7k1S0PKwgSIfAOy4L3ybb
BS8J6LKpEbmC1y84OYRJYB84sWMGemo7XxeJS2DMBMDIHgntSpjIF9yEMhYak1gz
1UyJQCz2dAbeb49VhRf7b6PHmk33zq2gH0jtb+meUr3eHlGAgfz2AyfObxzeDXHA
9Roo9AozZHr8bm5JrHfhPhS8/EILvvOzJSbAMl1Me6XQbRBrHymTsKCqfWoh3cw5
NOAOIKZr61ZtGI65s25Dau63vORsEVqy7D50rNH95R6Haenc+qgmlTU6ELXoejrB
2pS/xbGMlKt3daZn4vTrOdHUXoGTyA+dJfyMy6chp+nIsoh28Tp5zXLFaIxoGTaZ
Zom/6+YdTkgycFxU+xBopXoR2K2JGlNFraMyOhVzCv4lpsYN5igscT8mHmNXBQoF
c6ZfwN1gHhQg2l+Pc7HTTZYBSzW4UJDFiMUXkKtgkhq208pvYNW9lGSK1jU+psoT
5CFXPHivzvdHsjy8y5eJnKRSXvFY9HNpC+ifJZYAB8urUKLnkJ6f2mepbN+ZXH86
taT0mqphyYBBoeAEV5zPsAufwZAMgltpay+YdQlOMaOAYqn5eMRwz9XIUlBBj+ZW
YNWxfL5F4jRKnasjD4ydjBzE/UkZapGspH5DsV5v4pbz1MyUHNNBvfMoRLdiAy3F
MI+qx2z1gaBKSaqwrB6j9Pu8q3utqBx6HUtZdc/jadj0DkPQQl8PfUlpJb5J7pob
W/HzQaj2Eupb6DrzlB7Qyjf+59CjySHtD+4tI1AYVYfu1DfkX/7n1LaYZd4j1b8K
9vtqRhpgtH64QRvi6DRCpqFxffM03XCFDADizbjMIeaHEUZ+viy0RrXL0Lm7jgeE
qSaEXsUS10aRxbU4ZQMpapn6bb62mQEWPKnzPYrI3lJWv0Lh7Im9naFVcyIMp6j4
uU736HWGSxW5sSqtl9X6yuxKu+6WvKYFiedL2JcriCQ7HDJHiLrhq4W7mjejjbhl
LmAJRJZy07iJ9BpT+F3rgAjXsX8Ii2VeT3plPp+VbirNP59ZzzOg5z9KHxvxymzi
07N3SyXbstw3q4sf1OxYQLUSBlGxztFW/18iTzcv+EWLNXWo4rXdGoCewRXyKZJH
uCehOgIPhxZfFcPKTOhr+nyCS6Wa6l2hYen0Ee1O6O4w+dSP/yD15cO24YV/a/lq
jWSxaV/d3fqqyhJZC8e+QJuPCX4ouypbF7C/y4PuENvTwmgCs7k4L8OXq/xbS/qU
bICopiMtkRv8vKHioyiVXpffKHTgu1YFb+sKhEWS/JoXrBjKe7Im58nAgjn5HezE
Xp6dN5IRv2g5LQKtG0aP8zrgCNeEAkp3SbdQdrmYcg74k1GQWkwNYnG57e59YLn4
U1hnJxZx/l6Z8W38ZTFuy53HApM28uGI7ZktTfUd12MJiRjapXy/hqRL7Ik7Et2S
1/veY076MR5oV26fYWCDYvfZrM7P/Cakhy7ew8VEWsVHc9de2t3meuwKXXF5peWA
oGYqH3DNfOgaQ53FUyVtzrw6pxeatsZsIu6b3Tg3HHfUSwjjCHL/orTdmFeSvhtb
Iiwcu0BW3TCHvbqh5f3Lg/i5XE2H77i41BaKyvA1eAc/hwpEPmZMkg5rJOSM+oKg
qdNovauKUN6dExOeeWR6IvKp6ols131m4jcjvr/J6eAkqWzQd1XllAPiIz9fcB0t
hkG/6zRS6Vj4en8uvFCVfUrWjbWwEJFmLfhM7WeMq/dhxAFTb1CBucuOq7QGGMAn
GxUVj3dPPs1btd/75ew08LN1qiNpy2D9BIzGX4x5P26RI6Ej831gJWMzmJ449d5M
6pxrwBb76OQlU8ymDEX5GvjqpxH9bBqkCYoRSmMF/LehK0HbuZzL4ZzOc41Fhxah
bi0SWMeGd33pxKeBBEpx3PwF0XAiFl1Tz5vkrbKnebyqQou3++A1UkcyCsn6Fudd
fPQA40SWmnb5n0R4krrdq/rAL02DhH4v7pzNJeuhTGWgGsC7RDDUwNE8J2HhHb90
Qn0sl9cZWmweB1nPSKvLCYH1QdhCHYAqXnSC6/ExbtJfUsyDAQZ3RaIioR4a6uhW
FW8hN8Kj4Moe63dNmONO50SdToEY/32toSok5Gaph0Nkb5jrP3nD19yZL8OfhNXR
kebyZ+8WOKiOaLUzisty6ItpZ9Xx7g+joaN1tdSDMpo8yCHdcTBJWj6rkM+hdeM6
C6trBOTtfycMtzFUCWiFI+r+oqMdtLg0OCE+ipFKPJG2uxE5rHJbrfKpXITGtmWQ
Gj7nbk/ubnpShcSIZ+CC0/xHTOh0ed7W4dnyeeIc86UUSKG1i5NpRu8agFrcbF03
mIKP7KNRuQcWsdLvA8OiHw8GEoed7E5G5ld7cCM7MQcxpoYCsEeNtD3GVEtuoj2h
jvqTXuOZgSyRUH8TfsmnyeVB6SNDmmJOB+WfVTWA8uGS0qhovoEsRIdCdsf9uyuJ
R/ezYkICZFhC42Yil6CfU71OX68y5rB1VEcQNANJBM1mR4V2EFRzkqFBHQyXr4VY
Nb9aHhxyjxyMR1dk4FPRs19B8UghcfzcSBxg76BjFREm5oecJse6SPtCE4+R9JLx
OFZbrTThY8oQDrboA/lVeNaldrT8Ut/rj9svTD3D1A7HGVzzrZKQtaYMnYDiX9TY
Eo1A7MQr+BMuqLJjRmJsAqE6rTB2xCzpiw/CoqMvobEj1EwoEXQkN9XXLD/LOUQn
SN8FL1q3jZM8xPZA4GEv3YR+zqieGY+Z0Whv1XnOTuwqb7ojAySvt+oSlRJ4y4eH
lmMxFBboAquQZ4Oipj+8VnKkxrrXLsf9//cPjIBITCV7pYzP4MQ+Pl8HS8hAIr8L
r1x8b28cjIHrpQQLPiDaXG1ZOfWV+FsSFSELPkx5SPHqQMWOAGK1yAFSOOSFi23v
oasEe8WqFS8jY2g/KAUHZOAmqaKzx1xFflrBSnqtxuPg1l9KAfVeqL/Twdmds4Jv
vT9GIjkaq9Nqf/NoRsYIZMJxOUTh3Z9gwBQCbkPQxRHjnZwxU6gTLKYtfJ2HV9kw
St4X92N449eUjUhd7T6/ZJ6+ot4s6kt78kWyGi7YGH3FfcqBfUlOC1RKOe4a5bvK
ZstlFgbfnLsqbZegwKhcZtoGfOJoUJvye+TExeXxEGQ69GBrRrxztVn7dP4lnB9W
XwYiaTTP/AvE0SuY0wGrGDxoDpXo6ZimvWJJ3lnz2dKJeYYf+YjX0p10JqyGBV9f
nT1krygAoiFj1a8B/Aqy1bPlGDjW8lqHCDK94x9e9T8kgKeDSIcz1fqMzikG3Dee
B1b263DAngzcXXNiK6B1sR/tfjTNjWvloyR8EQxnQJfQX+UT0Juha74vkbdKo0w5
RjRSW/Xa+s5jbSp7NA+0hP5N4j0G1UrtEQ5fmvOhgZBSEHjl+lJ/2Y1MxAsd5Cm5
OsP7LeZJyHnPTvXZoD2FsZj9EL72JSEP+zVzSX65j5YvEdl3DZZVrhulvSn5AOXv
VwzonmolgfhsVKVsTeuXogNqZuKQq+CXMHuABslxX9rMrATdXdzpqvuoFQspYb4g
DzMiw/ijypuyf9AGCn5i1+eufXlu52b8E9DMrMrVbtThrUS4IodFmUPOy1atijhl
mx9AWxQmrAq9vO6WX0jqNqei8kklRr8GVtoYrjGxGElJIdIB2AsfYqiGHzBaOBDi
0SCpA6MVtU53VbgwbyE3Zo4WE8RJuHAYgL9jmlWXHwXLYr0ChEeFh+EPtHmfhZr3
uYfR7AxN1JA6OYovENR0CkIv2MfSNv2ZX7y+DCxLL+hBPHlBfy/YUZOcD9RNPDdz
YBRwqvKK1noqojRgrt8SwJ6R6IuXSTq3TiUbtnRSHWQwEe2k0KS1O2NAep3ONWbM
kXMEaKT0Q4viSziYsow5M2kdvm3jwrUgXaYqHQytz5BBkmQbyLFkFkPvLuBEXI8C
bAvbmmXwlCUxFXPd6SgSEeLuAMVdkqc6hd4wVrGGS5NSUESAYFkzxbx8OWmAYiXx
F14lDI/KTlLA1IL10X9KcrJHH/NsJdbtWjC1pdHGMig26+Aq7RH7I2WetWTTmHYC
I2khhJG5iH9RO9yG0df+IKLEiwPDisN6nMIk3NmC7nLyRdJGiKBiawjyCs7Pn4j9
7W54Z3blvGnWPya+R7AodYgfS864UHm2w+VyX/vxs0nzLuQqSS5m8p+UbH6NDKH+
KpypRuhOm7uk4X5t4OuO7NbTdBk9V4J7+DuY+Qecr6Z5jWgsh8ZQVEBex0QcFLU0
/mIZcRDlaeM9h4xmQUXqQwI2yiMk/2HjEMt8wZozaHcj2ewycBm75DZNDoXrEskh
F8ZUHAX7sHKwXJ2Jh06Zdb3cyNEWM9F2tIDWLzeTqjrCtmkyM4ZbomXEuByI1Mk6
byLtqyEZ2UCbMRGqHpyrFgwdZ/43XNp8EkJ95p6w+8CVAMbmdVa2KgwtcdEcdN7v
B9pESHyroUJXkjINvC+ZKiWzPQgBDeWToQfnPne8R0D8sAOiaZYkPk+6Uvgfy2/E
c+oxpDdVPfK7VY7ddX3V/kCIprLuMk3Hpx6AgzC+nFB/TP92sOhl+bmSFVj5lpCr
E3u4EiNmzMZ49bkHSamBT846HRlnJB8ttL6O/90X9Za7hAkLX29heWlfuz8tKXMT
Kdv42LMTRLzpeU8Fh63lSKi1EVtkYSl94KQsD2rVLD4VbABGNYu6UuqogtzhwmL1
fAgG1R2fQ2oAAU7UjCpV8ZTlEkLIZgUPrUM0WOkJlyxKzKgkyM7LQxQOwRBSAqif
sXLnBt5abHeZlmZU/DgIY+cWBpKWXm9XSNg33vBiB1idv5AUhspYp7NT8NmLg3du
dpd+sQjrob+lfm/ZLV3k41bhrBzDfHQVeXasx8oIW7xGUl+zh+QRFpC7dtMjUBXK
/sWN9tkqmCfwwxPM0DdKWmJZwuq5UCY0tPR6MsRAlenP2aq4KLqfcc2JOF3Vofw6
NJG2YYLgLOut+8wN7ZeOSqPiXbwEWYGYL8X3Bsjrc5lD1U452FdH2k2XMjVrMf5X
hgyO0a62LNQ8CFBD8Z4xerBtJ6G2aBpsFDcmN8wbDjAiAVgJX4+NQhq867B62sWs
eLjNgVlNgENbKudxZ118X1tHBvr9gXox+fc1+OAlK19layC05PA0s7P4rokJUv1a
DFFA1zzXBBJPkSRVPfPlzIfyzsJIb96UbnEDc82G108ciFodo8I4m8o2ogXCjWwj
o67mUX+gLV8rgb8GYY3ProJnkscind4CxDRp4NMtURnjRgVgpH088aYwdb143kR1
i3XzPtlRzJ/uTUQuyCvJ+P0FodAU/TtJAtlRpdFdYQOtnI4oqLdQ91eocVuyHkoC
lyzvPuv6ecPrv6uMVo22/ed+55ByDAPmT5fnWLJ/wK32gYQE0tjonv9g49oaPN+d
ba1WwkeJx4Ya7Czo+gZnewBqTSlrmN5mfGESpo6mozoYUOEZ5YmVA5rw8UiOQP+k
RLFoCMYdGa2dVTwrJ1jyfwUI1qgLrGiUU2TSChwAnkX5g5qO4FLZI8kK6FGNCafV
6wG9/hUWazDnQYKOdOiNteE7JTjHHIhoy7eI48WN87/Qk7NYfNWZhFuqcjHeZsiQ
8ADcODp6CVePr0bifMsvv+6rJQNAJSoTg8dQFnUfuR/bqDeV0c6PZpZkfdvziv5J
DnWAVFVDYm7Dlzi4ybAn2lCddjzEdvb7tLROeWm6IlEHeIcVIRSm8mvGmP1MzZZb
ulehGjkVaNJgMonELn5eJLfZjZi1KbRAQhOkLfbiqw6DnqBkzN9gnYiPyXOXC520
PnBknKLVuF/anJUyteX3CBTbb5UFHzFmU+lxiYaplfee6aUyUyXjvh7sAxhKtYjh
DggssswbNDc5z1mmTTx2ZmgG6jxNdi6iOwsLNaaWlsLAevF2LA8CsL+zjZaKw6m7
2wD2RZVBRoaFFQ9WgTCvCy7gaVwMbTv7ovkYyMvpQ6poQIe4u8E1EylQCt20vIX/
GKRIgC4JPTK+o1UJNHehOnZO5Q1EQyzjMP6nyExdzn/uWLYoaoHvRvQelb66PkNS
S6LsB1NA1ujnBpTfUkPHR+n9c8LLMiEeLtSyUcTi3qzKf4Vlp4UuqjW9J2GUYRjZ
ZSJLD59DANlO5bcOXINT93m9fAU+i9X3SFZsM6RpuavRdpng6YIhhpdgOOBFZwNw
WoVQ2xHMbuSWCstJOycX0la0WP315eO3TpU7l0yrf1KnqYiuCLz/uy73T4+3Rc4S
2TP8WegXHl5LWUN6q7P94q5oq7s1E8LPVnfv9zD+ss16F5BtrfNoDByRROQu02t5
OY7G0ssCLz/8JMo7RT8bQR4ZxHKJC1NI+toLjjwSUxPSGQegyuXfmgAeCOepRc+O
6TZQD/hw61tH+8yEE4CTqPIvC6b2R4l0uO9fuZwr5fXzzDiIR1KiUue1HCR9i7Hk
avB2S8VW34sxkOTmlRTKp79KGW2V9VDZVhFHewjNCledre9YCvOUjxojqnlNohyQ
n/VndfcN8TBeMqzFFpDlqI9cl0OcAXaa9FAFG3tqOBz/jM+UGWA31rmUNOvwRGYp
l36KglGTmZGQAQUsJ/uKVKU/GaZdCOJ5ObLllNjaDnuADP+gq3rVu+p6jWwmyxiH
PkjMQLpgEiTXhqGHM5mHtaJgStVSIDVlVaPH0v9G47zCPvelG1JlBcHnE/G0cgWV
IfoRLG4vHEmS0HnVT7x/64HWmYiqDHn2vpw86l6indsk7NP1RtOa+2kFTB7ylrvh
RZ1ymxz+vrrP7yNr6BKBj8xpT9whzQRniaG+Ur8Fn6rH3oLYE5oSR+ezJbfgU+mm
xB1HX8N3pvvW8i30b6YCkVweWPfwPc803n6Wn0Srj7E4EXH0hGfn70IWph35eQsO
ceZvdCbvEX+yoz0vIOvBgmMDQtq9GOJ95B+fJYA900XLvbxnssDtDRCqEFjnBV+V
qjr56TR1gANKS0TpaO5Ly/i0dpA+YeLPawc/sCy+ijHfZpfC6GPzsT8K06FoiVoA
ja4lTjUu9dbMMvV6t2RxOY1n+gHzPsOeF1CtRmHY2DE5xQuELRRNf0A+uV08rqKK
J6QAdW3SYSZvOXgpSAM9WsZo5hbTHm38mae4dKs0VtaI50DSpyh6+776cBZq5QdR
HDBVTzT2HJ+WDUPPXxqQLe5fPSstb0lXsKS+nxqC0ui7Hf+9qcFX4hFTCQDjAWpX
wq9uAW6CaPZERAiAa597Ad09lc72m1g8qH7iNQd2wndYNievoGRRFFCvItkzJ6DK
kwT0Gf0e+bvRwpiWMyfM9/Q3l8Frk3c1pUF9xdvMCIl/cLVhFIMaJK6jWznwtXLw
ftRdIc4WXLhRcWLD8nsgCEZqBYIhAN7h3//0uzdxo+xdDqtctddQLDGyO/dqKEKv
qzSiOf74NIko3KuH2fCmFeSOGpox/4F56PoCkICgcjc9RNiJYGUDLNSlN4el/6f/
PcMLl6eVSaAXdk8AdDqk0NufwJeTWNBrYJoUbZXsfbxEHt8QDUrfLwmpzN5Zdf+U
lI+sBe2NrjdU8bmE5IOXB26NjdQiYmmr2cSSjHxosmiRJ7ysnEbUT0Su8428OUTB
mB/djBOvJEMj60kvjXJwy2P/OWFTR0CWx6euV/hNXzR3ZIl+4S64c3SLEZmUXoUa
bP267JqveGqZIJWBepwNQUjOhDgRvLXdz5SN57pJVLjsbjEkKfOTrQ5ZVq3XiCCT
UADyDoEUZ8TEAGn81ALnUnkwKAJeamwbzrr7Js14Hdm/geQAloOGmFxLVJq06Pzi
gHo2/FOKzFY+W+mhtvQ0FZAXkwWh+x1SxuhgkOAUKL2RTsaK/vZeh1VEqZJXaLCH
s7IDF1uS7H3WxEphFv+x6Wy+C+s+nxJG5aYHdaPyqalgn60khUT/LKN8WTrorkkY
bg9Wn/rih8N4IKgSLwq2XAM9m+wnLXZ+B64Vfp+I8duNjE2J45J7v2g8aLHCtN7K
ZuMd8Iu8wvqobBdDH82R8SGph6ZQfyDZAjfMJGf2d3O6oT/B0tGscEkOKTyzCUrI
QXI0pHfYd3xNSA30i0/nG5V2Dwu1qZkHfAeNNRfFcLD90Ev9HRKAoG8VcEjqaxzI
9VbB2Zm2WMgrg+QvpJjQDbAt8tIOWcEpTL7qyyvC2IcfAhU3pjGl/3QONyL+m/cB
fwSlO4CGnmTxXl2TPWthUlv7QI/Z5yHnqF5UGw5JqhppEBFmU4HFs8S7XQ12O8Uw
KWbFSzgAphJTlHnHyu2bNFHq0wN7IKff115abRKXIYiZC65PtfDAiowlZvYTKnVr
EFzOqdMorp5yXDs3D+BkJPd+J04t3O5uXeGK0D/9Zx79HaPx80djZ+hRY2p6AaGD
kJdnZI+d5iG9FfFWy/Z7gxHZ/+EUvwDJaDZ+E2R8XCfVnVQamTLxYjQCxLoEybl0
1u2oFrH4pCGV/I8/4Z+EBjHpWRk0SohLRonyS+DRxFxlm8TVvf9WxFRZtb9R8UNx
NmnvteZxXz0pPxO8bRVsGKK6XikWYxGz5nZOTQJjEzXZpilGgFmS+bXsO1lNraom
guvAQmjGsqB2WDINUI4bqtHJZkvS/l/NqAz0Um1rS+CQGrpJHw7Plfwd19gMK+EA
RH2lngBQydCmB3alxqW+yjM9UdPmeku+4ofc4RKw4eeXsg9TCuhM5IocriplG+5Z
78s6BZGB8ahS3blsngTGomU/aGftOEVULUvc3jMD199v23Nj2i1HASKZpq/5YZs1
/+pRMO9tpEPjsN+0dbafsmN/4PKaW7vGWlhG+rAIc3D8VS95bHKzSTPYpEL/zPpe
nGo3N6sNYdG27zOwiAa/aHeUu8pki93HYf1rKWQ1fgR/P1X1TDPWmqT2qH+iIiw+
ui30iEOti0ccNnzaoR+3sEbAUTeTNPBJKIrhYvRFPwY6V2FEkrvdpB3alX3DPld4
f3eTl72AXZTtmPURu8XG78QIBvGBObAPihfPS104GPXxOvMqgRSIH4g4W92iYv6l
5snMkq72TcASkEj0hCk9s5d49iZrAELrQrPYVOe+UBWQcWEf1L0y7N8HsycYMGWa
Pbd1+X0jc1h31jCK8mhYDY7sLRtJ7vlUvsEOU1npKCbHF57thsZVxC9Og1HUQSTu
tcgY3/WGJxczdZUt7P2FsylaKE4VhFxqzZlqGleNOCzV9fWO65ZLsvwj855A1wfF
qMZ406mxaOMq/ca2oGA2YjECzSJOtgvIFmJYWZyjPPofamPU9kvVd8F37rvV14Wq
aQyTwaocWyP5BfuOogXlORwT4ZCKT1KQAD3AeG5uhG7NmdL7auKxMY8xDAA94tcy
JzkIlMuwq3muoFR647Hr3qYIZHEl4FVdG2kvQjIXGc5zM/eM68jgn4dyCHkCrg9U
0QW4ojKAWiZSJ/ezCYuXN4huIICc5lj5y11+kifyKtwNuS1HR1ppt5ZfF5mvydSs
0lCLkitty4dnf75AzMvacrTCilLWHPluCe7M8iycbfngj5V222ihfR5fhnOCBJSo
PjlNds1CUuv6vGTYK/P9eAJj240Ose+bY8IJnG6FQg5i0d1q3oIFA1PUFfvCWN18
Ly0mwJtpT5vybBTqjqQ+mk3fai6em4cTgtmR3fEhhl0FoNP3FO4o0ZFelDDOvCV+
DgedZmatNDMswt6BcJQKKS45Qbho25kXwPlkmZ4019pV8otZmIPmpEmR5zdhqWJO
Am6lvVjIAwu6SOrVo+nFM1DI+jXBZu1McShXaKp1VNxOj6lecwgvHDlrRHDAxUnz
uakwsx+hij6/xmkLXp/ldxwyn3EkWvfi7eFM1roGD4HVThYgyf+iGd/msaTmQEpV
b2zCi3zy2fmndLvhe31F314sl4PcUB2sFl421QokwyBr+R6wVhdpij6vpCAUKVE5
nkedvlzhCXkkfDKdoEQo4cmkoC9z8l4IWnqb0xrn30awZL0JlC7hJm6yT624+2bX
qugUt3c9xeeljVqrJUG13pZZGJd4MY7sdIzE/6ZDyt2xBuyWNdbGVjp6Nu6Yy9/1
J10jKgh8+hUhQgxTHePQd1yMgAYKMiszvSGk5UDoh17xAiqf3tMwsBMSyeJT6DGf
roGR2tagFYvkAM25vo4jUU0SIO32q09USZbDU3RKrdkXDr1Xlf2fScdO9QNno5lG
hnSDFvY1BeL+LsTwENyfcH7iLxRrj+W+GiRSY78OjuEX81gSKDU4owMKOboDw+y0
02tyYY4pYomlHeqZFhkjmL2TqXb+itXozy3q10fuwVyb53zaHKwDU1EVFhgghhup
fjQBj53bBySz3IgLYGCRVB7vOarwFHbJKxBAsSMO3XbypynbZg7c+QFpm/G43T/A
1AQM+0/CKfAQotpKqju679G9fCFkOs5Vi6GV4am5JM4Ilp9UIpe8F8UZyVjEg0ow
a/E2ohSGASN4DcmXVz3MmkqKG2i4ikaU777c+QLaY+GPOB/OOzYt33BcaMeFgc1d
Zj+qoGGtoYNe/WhEO1qbLldvBhG0Ga9xL/4blVbRryv1ytq+UITH4NAh0qXHyoAJ
bX8z075SKkZS3oESYhA1ZfHKNzz2PZ/Uu/By2avIy08RJJK10axp2POEVSU9l/em
ht9S8leEKFHCnZyYVG99j8dZFyc6meJ9QAYUdGGAYiaY+PjU7D1tbP77N13JrmYj
h+s5j1RL+vLWClEdZFRtcgAIrpf8bHXOMnRTUnsIwHIQyiYE7jZSzmQUxsuxn3o6
6/QlZH8wd50PNgDjeuUbgn6K2Fs3z+YrsqoXPHBzZFVzfRtQEiHPuMlIjr6gpxf7
CQMnhE5YovgQKX2GZvYjQ5DOJRUlL691Wz1wQW4Hp5J20AOJaFx653uiieHtmoh6
NaNGKNsmSt22RujRJ0Y32Xb08LR/ONv9u6Mtp5LUPp2fEFKC2MuN0NSnOWdB2StI
iJSbYCywKBwN7TRG08QBm+9RmHdJfJYgc2OxUX76/OdNFqSGysTmohETWHQgoy6g
xsElQjJjWdulfV7tO2RioHcOwv6psJtC7Fr3rJOzJ3DnWqL4W3Z65312h2nsP8yi
9qQNLF7uEONMTZ7OZOglWpG6msp6IE5dnoYLlUivAzhwfCh4Jl+rvk0E9xKocoM/
g/GDYjDc5vfrqqDZRcilxksO8SLIP1JNvuHydUsKbqTNcoOfclOCOdvD14sD5ouF
o4n5iKgLqgdtSFigQs7PgujzIS/GyohAUFKZW7nZTklvrPIuU/OMjSckR1fdK7ff
tsY1B0tzLAOv31R22PRqGZm62NBgTR39xLXHBbC4jw79HMK8SEG98JLAuSUK+o4R
Q7XFs0liaWNDY5POIj/7FkMbhdatuiMciYx8qY7nPWtN7R2Ma3LVjI5ZQuWhfjt0
G1qZfOLsXjg36g1ocR6IHpAsGEli6bh2ZHpUtmpLasOh1NZu827OwQckevfS+93J
A0+fjkclbczrdHf0AATTQPn5E1qIT+TvfnyeW7tnQRBR6XIl2/JGHrhrb5VhKMRL
FvRgw4KHf2GjhlxKj4eNIZ6IfNgNOvIBipdH5Ei0PCn6+NA7RnUoWjnuFtj7csir
1S4lt3uxDmLECYyP/Ne5sgkcCqDIHGhOeOFNm3nyAXdiPgCk1WSDE3qmocNY2+d8
K0EHeLxOrX17VefBFKpw873wOv1JVseNuaWwb59gVQv5kOp+oxka1FnhmxyGalf4
vkQZnZzoCugurgRSwkArgltStPq0XPdD3xraO7fVgH5ExaDN5z+FM6IOHT//pnmi
CFf6rmbl0iyOEZupRc5OZNnlm1nCK6abl4QoUfPw4QVEVq5SrBG0Vk5NUqNm2Muh
vHyv3FoYFCffVMXlbiYkz+OH4K3gBXf731wqGtPtO5XrMcMN7WRVuX8W9ftCLVsv
TenRG++Ki3+3OsgH0Vd05YEdHN000k/zuLTeRxhAmCV8SSDn2dMR2mQM8zEmlWZz
giatAcDwLvb7YsQzb0IBkhfxdXb+qCYILxmpykUjAmtdlpSiVmkwULz3vWOIYvrx
wljdxo5kZgVjSXHiHfQVESaBJXKoO3bDzahbybd1gr5poyM0oMNF+lN7ctRS8dxO
U7ahedK1IULyhtX1Pj8Y/bExqBSIf0ftscrc6V29sfA56QortvATkUnD0wwDKa0D
3fKzTWqRuQRQW3l9v4fMvIxjGhPyh7gOOyQujjvl8p0VTSllNElaiOLn819rKT7W
rCwmNjxnVm8bJasqe/cEptFy+P/2zW19P7OZtaZm/EKQIE7aVxgGSkNgvausM5xZ
ASUD2NxyRfU/3ALhgIm1Laxtv84Vlul8b3UXhZFVOtoQe6FOLrLQiCE5n0KtXLMA
jN+PW/gJDJ2lB2KtGQ7OdY5B3RkYMyMOCB9PyaJ1l7k1IdM6uMMgrThq9GxoXRof
Q9cquoE2fWPm/Hlv6CiLj1p1ZdAMzDvpR2Ry3aFSOJQ5XKukD/hGxH8p8xb/PgPX
ckl3Ue79hQqrm8RK6mGdNiiO/HZ2R1iHVYdaF2/P4AY5IuAOcGc9hHGlPoI8GrY9
KsmE3Dzo6BMPJzgPEcTGHxcK5U3SUA0YEw3ctEjvCSQEJKlNvwKEwbHWN/gCvRuv
Mx0UKj5W5uStVzi5q16oDvgq4AfvEhTWq0UDa79ElbuQvsnLpnA7iTmTF7roLYig
kLBJvp0w+mx3qDNJVFxHoBzi+SZ2wyJuHqaa3DjNF5RrMMe9J4OpcGrmUGKn1U8F
jADZKvy+Ro3n8bDS+COY4SXGWs6tccXo2TUtPB4HO6KVEUg0DF8Sdg09aY7FCqsa
prxyfHy09jrHIPoq2kJew5t7xKwBLrtE9d+n7BxITpdCXcXqlPT0ky7EhU5eWi4b
W6l42mion4Rn3qx3plJfaeTs0kHzEGIxmUH5u6ldr5TVxfO2ldfgoGTA3OyWImqG
yWOeq/QyTBIL1PGz0UG3NDveSDf6KcI1gr5FTQC+sMfU+l8lbpDaO6B5NCJsINu1
63r5t5xNiWM0nEV91ReABHO1s5RJxO/81bedwDO3oj68JRH0yL32dvjLXeTGOaPZ
e0caY3WR1SqxQ+qUELaTSMEljbpO5XnV4GfmToZDjIhKnXusKUkWvcn3NEYMArHH
BjtpMu359wz/h8hjYrekLHvkJ3Hkn8XPIBBNkqhzdyfSDjpOePcS5Rjc4E5VosD3
DaG/T5zcchkkLkXNIwR7SzbZ4zCN9CU121MV/vzwFoxNqa7tEv9UBWr7rwNpcK9p
6K5t9vuOk49J7RrqfpyKOXZPeOHFnswNpU6Zkxd890+byU+QxcARh9q+wkfFazmj
J6PLYTW7u+aOPbBGfey79ioIzgo7s8FhaVzOelty9o5XTi3pkAcXE4ublexDhib+
knXu4fbP3Lx5ge8XKJweINPqTaBdFjhtmOhQkGmsae2NlLNeGEY71g0CVtndaK7b
/NjJiz+69WAMtesdJ/n519b9EeYftAvVBmvgCeCQnPpxVaPauC8+VCvl4BZ9kLp/
z0mLChIiIjdOJ0q3cbBlfdQqcVNEhMNTOC/0gFMgnN0q+6GolVzQSdNzwy1Ird/Y
6k0Hi4DrUmpFs56+K3gKkXZzLbzu8ffV8potlqjC3dp/drHzH3DDUWlNOlJNv2yy
xijoGPtKQT8poYLM/9Jgv4hwava37hnCnaswbSjnchO74ioIwLrbweWL8049iYy7
N8yrHui9QvLJcgyNdNr80DjGgDVAjCYy7SR2tNuLbqf/L1iAfAsBWnTv1Zm51zE5
qjlROt6/0Ib9O+L5q/r7fYs910+AmQweO3HzCcclb3NiuZ2UXZvFdDhKLZXaYbp0
/qJaaWxbbTKRUVHV3CtvN1mRu4W5gYW8zvasYaUJAGmX2sMjcdmfU34t2IjvNDcr
f3zucLJgVgIo9vyJofxm+kQqIOiRDqubuiMcbHE0IcoyBiWUqhkkJ2eig8Sa/A0c
z/zmNzkc9BmFU2pCq1mUa8CHuIsiFx26g/fDLf2BE7v/86sngm3hutOxAZguBOnH
bXoGA6DI73vrhRYaMBQ0oUS4hAsomJ2ilHrLe+rmtfxRMavAAdl06OdkBMuRFD1P
lJ1Bd0BIsgGTT/FQApdNbKKGuvAa7m3JR1aSzIkKcO3BvCTyB+2MhgGeAOwXXFdM
JdGlmGSqn7y5haci1cZWjvEt+CsBy8dIPuvf+B02RZMz8G6Lhf5vq4JGa5766Rso
TGfvgwYibfRdxAbCh/Kh+iDWHEgL1Tt9sJIsyUYPw5gHJo4JlMkZvEkgnyG5ddb8
1mEdVydwci93DAUxANaJ8yI9c71C2jHlxBxUext9gqmYDWuClqMxAc7b2RkApaNy
fsUhL05KysO1qGYQkcFqSbuEKxLRvk/KYEcfGtRD7/k2z/HjZrepFJ+QwSv1esix
q2tJ7B9DSxyA+wieeevevKsxZi9BHRDsAtJnoLOciCux8jFy/OcushfyFW/jjpfq
jfu6cONf+NOmDTsIRqLmSMHKfPPkKmeFeANknHXOI0icqyY4HJOLk8/MRR91rr6P
8bGbq7wPRVlValti6KrpirkXdg9gaaZTkWNRSPWF6yeGeIX9b/xY5TPKA75EW7Nz
HQzJfI1lcQ1RzCiBjKotV7UUkWOYMi2rwqos5FWFESB7w/JQTPCzrMrCcDdaOKtx
bH95TLyKRvdYm6AdodaFzOA3YKaqdnABfGfa/rtX1qjmb0OpEJX9geKeyCYJpt1H
Mht8bGDF0FE5exVFB3dU2MJfs4q+bLDPqimcLyiXvpIkluN+d7PzQ8HxA8FWbtXG
Y+6ZHyUxcFLxlt2rXpsQs0m/09OtC3PI8gBIpVXgBpQLTB32abx/HYmvcmM7t0CS
DHb9bxNRVntn6jyCd0tYFlPiUy0umtRzHNWcIOH/761yj14BsQX89pPweMn7qXW5
7agQ5xd+mmZjTzOcto2LQqz5J42r4Vl6FyVNIeN+wkIOjnhOUV+474nHlr82hmNy
XyF781aI8NlGDS3rsCN88sg1sJNNigMwxOJCDSg5tXxz8FehGRpapL+scVzpHTAk
wpvLUmXIFI53Qpty8gY/3nTk8iKmO3C8bGtHDDV+WKPIHGAlJ1kLz0Vz7FxacXcT
JBh+51mwgswWdvlxN9uioJjO7X8BBBSBF2IlUAtqopAvtn54uezYq44Dl7pgD4EX
pS2Vv2p/0+4+w4Y4afF8jj5YSGi3ljfNvMmfo0znnE1DW+iSownn9zCWG7bvvhr4
O25WyoYevOx+FWL/YjLcy2MnOxSn+sNw2Jq5S4FekWfWPSjkK+nzMn5GIx3JOinq
hNlT7jR8H38P5m7r7aC3S4uwkRsTn/5Yk3AhfzbezYA+NocxdrHI334q3gNe8OZH
ZDxMrGm1lt9p8SvMcfIoyL/uTSUN/0FSDMZKI4/+Z/DLxUB63ajgZM8xam6r6jP+
O4PRlwNLsGHAYq9iYnFbnuzFpLwH5SEe9M78fuEs/PgKZgTJ3Rt8FLqkLl2vVR6e
rogcDKaPrNUoP+rJrFRz8s0uROPB5nroeeAhgDcCjQ2NzC3ShNAkfgrfnzUq6q9+
xNj2wR9qu2ZwSpxqKTtoZ3KiS24AK5n38tYp1LbgDlWAjIy82GPTbN8TIaxRVtX8
QifrUDBGskZzDuEMXTkVir0D495JWqSEwoTkXUeilkhmae7PdGGybqUIO9I3RwE4
GpzA27UubDq+8xISZ5EZupnufg+LCWv22LZsLmVtT0/efO82GMPGXV6b07xa5BU1
dFqUaFL8UgNvpPey0BK90ZyxUV7AtEwcyTYq4BlAYq2Z/V7575XCvWu2AA+Alpa6
qXjKZ9xRLZCGcGLoR5XPqT2Ru1ExbaulIZNZt3mP40pr5fu67NOIt5KKQnPDmnbS
+R0ns1fs2HNordEErGjS2LAGMOQyUZUziIJlWvq+X+CEPYrA6Qp+r2oDCDNHbCKd
+uIrVibYAkqB808NwAB6SxsVU1mfoD3TRCfGCXLTnxxDG5WCMEqH8Jpqa0bxr1L0
94HwFMI8yn+t+f16wjIU5tLCcZJhecQkWra8FRWDo6oOz4XtxIimeraqEusPa9dd
QNQV44j4uFYdKKbJ6ETmez0o1O2x8laZzPG46JL81BwmuUdfBABHLgtt+9idU7dP
61atP9OotM+zW78PbnS3WcZe54yfQ5d+5uG+luE80mZpqkIfrrCEMYKGJKF0sA45
wUHNPdKpilxk+V7FWYCDpNrTTvdFHwKTRtazb4114i2EIWpjJzzoCPoYzrvTeNVU
igq32dVPKOXIZbKNYlMieZDOxoNyWcF5t7Hki/zX5s6XaaWLkdZK3vho3+otTK8S
WvXPc1NhaU9tMzFSKUj5Qj1Tf5RO6f5wstIKiQUe2IZeZvoT5gkyaoy8QKPVdfQ6
stUCLth9ToYP+GGozXemTv88428mYGQXzsUht2TORsXJegTrJGjJXbPMFWCHFgFC
Nuuo5cvHl10osHVn+xSksbcVgAhcRWNq0qLKJv//kca86DduT+WNRjPamDTBvLfe
TYaL8//2Vngv8NuwAQ+z0Wl16LZcuj0uzsz8H/122mVWaIw3OKUbAwnv/bGyhN12
bT8+Hv2d2RJRYHnM4oZqh4XnhfDl1/JRBBa1wTrhJcaN35jLAQhyqwhWpayZOd1I
Iv/AGckQOCbC8ZeBPDPvpXtLZ7vYHLuaGZn6MSBkD2BYzEaEg78p96aNdQHF5JCw
BiADYBMpQcSOlMxYeaU6CuAnGfbXFQIQTP40ql0PARdh/GLhAcaWlR2GZ2Tgy60J
FSYU9202tc5yCyAIHNJrMxGtZxubgvPceb2fMb0PZylcizSTo7h238Qj7W3lYBn0
WGrX99vQ1wUxwNXANUUeJG/i/avrmHmK60A+mv35M4qFCYJ4Qbq01nvj/Vzpztfg
Lmf8C0CdSYl1Ew4wpGsPpLEf4eE1X2m2il+Sq9LvapEl9ziRHPJaJ1jQI1XPOos4
vPb9XPtwZNtSJuxgU4OCm6o/9/pvRw3ikuvRKxiGYeAsx+KzQKEwXORwCYtW3kqt
alHWoUFdcLxG2m9hkANom9LRzKkwnt7mxp9JD9xF+W8KGv2V62poETsejTswDSto
YLAONhh509WoKgDRaEVP1AngvyRrE1Be1GEm9rgARDJ0ZtTCXuVQ3yECSVN8ctJD
D01QvEjwxwUn7vD+QQHywx8yTHfSq/wArDpzJtll8t5vrwr84+oXOjcijFo1SM9d
hjkz66nFT7eTjcxHbOf57suhkdxujEEulr1rZnw6CvQy8J9XpyUNP652HojhiXYz
09QYCwcWv7YFmjrwALAasWePmTT8GJ2D19d+oLQSXW2tihj+/6n4qUQtG8ybtJSa
bUelp05XWDNsYn/c/wPZcTsua6qtvMJJejDTCnSTfoSAjPTf8Ro1ZJ+69/Lcje2J
q9Ev4/1G5cN4rz56Pp/cq8P6p6qEKyajg1z02H0wO39pF8yRTjAnK0IbmMzomqh9
IwOuBqpswsdFxXA0kUe2WejZtc+/h1jTMzhC65QgQK5QY5sSauhBm9Oh5NWZ5vUk
nROPs/7rcUp/yS+t1y8fZhGCPkFu2hqwp95etCm+Unt/oprJ2XOB3SwIVCWCxyXx
EGRCcaeS+I56lt1A7FuI+ET5+AsnT+zxQYQupGinbEtUAJ/cHzT21hVqN+frZ87+
hBMhe0Tqxi5teRpYNKcWcy/L0Smg93dvB56XrxdHpU7/w0TmBMH8Z17aFLglTMOn
RbdVz+dDQacuo9eYPb7YkPbHB1Tzcn1THcR4aqaeAO8l5X9/s6XDtm9xwHOB1rpA
6wk67Y5+lQ/tcI1+fBcikersWTHfCZtWc/Kz34DLnL9G9pdLDAgm3BD6S2y4YyW5
OXwAVlRmm/7DDdLe+VQxUYkRlKKzcNZNkV3+K3yv8GokEIjUcsELFjOqESsdB10O
Ba9Ipl2zhHlkj6KKeLZlfgCaJEX1t/x81pamK2D1BxnoNv9guRk3feEzAJf1KUYz
+OSqnJA+KzbE0If2BLCNSXC1EROGA12CDkWCxkmHcF36BJfjCpIrKXEuN69/fE8m
MZZOEtG2e4H2Jk5aGAc+92+6jU/pEf1C90EqD3Otl2OzpLL7eZT8nY6MzMqfvQBb
G1Hz5NVKNRfyCpiCh5x2CkXyFQPVUNfEcltWGjAAl8unzpQPYmokO89kNQLiHFUY
hCzcADUlojPAwb7wMLQBK28237y51E3HXUeLapk6mob5ieweHYMMJ6U/7US5Uhqh
rdZBfbukaVNhrv7R2fZOaisbNJ8SkW4bm5apes15wRosXr/p2YPdfYIWm0TqbH7O
kPHU80hkMq3Bti3n48Z0diNVHUDaAaN4t838XY54welN8f3CDYtJzZc8TGcRAV3c
ZcCfdS3SkrqlinUyvL9Xt5rvFZDc2ECQaElpQ34IB3bIlwQoQtzFeOWk2FMLN/JI
wwrBjcChID0tMxuyFWpqfjAoqGz//o6jrv6S27VD9b+JP3IL1CXL4eWpdxpsvX0X
5il2p7IoSfK8TfJ1tsQBSaXijxQYHfrT5//hEdJyF76q/UMZ5GkOPNv8qUPSRj1l
z7qhHy3YemIm9kwKwlpwSBZIuSQM7Bd7qmMy3aVskUKVnoVxPE3QPocKQX22e49G
Qpyi6LSGSlghC0gAFXWSBn7QKW7UpZeTSekM0j1vpGMgZvsUenViNv9L+IIBzHas
1p6H8QbP020VTXaCc/4G86TK0HA03IKk4SgOliH08NTt4TCSRJopLJSGbnUwAse8
az4q5nwoktk8HT6vXRRd2f8Ts+/otqBalMG3x/RTbCd8K714NTbIS3etO+ULZjq+
+h5E8hfAuau93iTGfWSoZq0N3i1ALQZLG6yaevABoALP7sgn6mtXLLjbHAPBgvqQ
0nM8vPnYKx6Hg4NgsBTPQT7uVDW9e9AvsdRj6Is/pGjk4JXbM161Ix89eHfQKSxw
qj+8hOYqXWig6DDt7OjL+EQmhrKmHzqb4M6L70wEqpNfD5CxeSKHySNTUjshDlie
zpMV4ifswEo1uiiRsmn4boKWa099lTQ+ePg6+7LBk2aS4V42PM63Hqod022SQWMU
DpuNrT7h0+rtTGURn7qWO+QP0WVxsoix9rq+zs7o+7zniss5CDbobtmQ+rmY+OTA
3/U4TO8L+eR/2B8f07Wu9Low4CKwmUCGvj+rPl1ARbKVZmPt3/o2fQ+NkEa3uaoC
5grsHI1tbItFq3QIMh5Gldv6r8knc9pti+mrIrlWgFqM2s8j+Xzaz2ONB2J5JR9v
27n5F/0Gn9DEpXDVfnmDGHTr+t1bHXiBMV+hh4F1NSJl4mzsR0rk5uutSCxcakby
iO0n59jhJn1GwKykEoAwfoY2Mw0sMomdoxCa9c6YRhm1gE0gsixxB18aGynz66jb
FHLOn88q5e8YhvaANNcHYW8N0cBDv0Gc+6DRQ7BMs21/gVonufrCaGyQLxQcIJVP
3ZNnMkvC1asAtXtdsVqxqsuD9kuwMftp8/sSkmtOxYSWWAWdyZZfLz1jF/UjzLA0
IIZHpeBJOFgmGDDq0bDR5fiyNY4l0hH7cgVtOTkNi8enzNDjnkBIrlJ+kBm9UlMc
AsU4OYv3IR+Ll8Eu+5jgX9tN6IYCmESUGCGpav4JA3ev8Lf9eLr3SqMT8IbZtdcM
CpAeXM+3lHJrphLclA7oCrEWb8dMPNBgIJvK83c4URQViVq6L1Y9aS4HroLJOVl1
W8ZAFDAESEFS1TrR+SWLPmWy+VmVNDbkogQaxke+o9HSLp+XSHOgAxn/tqn/0DIX
PI6r+V/z+3g82Awf7BQKNyK0Y/jhVzwSfEwoe66doPMuptVbS+0RYznZTTIzmrFz
FhPxSyxrX4SKK8JU1eEt37PNAg/6984aktTkje1oxCYYRAkOaJZjgmfw2UO5HJp6
zDZb1XypbV0chGGU2dIOYgsQvsQ4f8dirQejR/kzeVr/7lnCJs9n4CYZOa9myz7g
G/ghuhriySy6BJtfcQ8EXWO731Ag2wpDylBRpLkD9Tp0x4wKo4xZJ4LjNQ2JDuzE
/rEeN8nsFmQ632MgyQzryvrCNO6XiENWni0w645BfzaRT4rRrVSJCNN8EkGcUlYQ
NkPwh2XzB3hvq7ZQ8IyoKAGkXiZRirLdsnMJVQz/95lwaWImhi/qtttUS21ZYCed
QX0yEUZdnGsNH/tCO1DdNHQzeoNuey+V5uDq4/fYhXbDhXCAaqHTT+6FHnyeC/CO
T4IG4gahWvvEMyY16+qwyreZXKY0Ggvhfq6BOMv9nu9fpI3OpRUCzu/FeceORCDp
pjZ8e5MXDxcvFGZlY9mU33spuuvNGQea98wSCXlOcKkaE+pfyZVhbl5/H+MbqtI9
y4kaoFolstmR4yPnznjRuP0hcOL/t5OwcxySKj0k6YJKDamvJlOw4zkDv9KBJNsT
V9D3k3svnZI7nt31bzvFiMmCPj1xCYU9g1IA7Zs5keYzoKWmkvpZmXyEJWRZa/LH
O7ndTvejurtVh4BVtcDaP5UJT+Oxbnv02BrZHHAydIQMsmqQ2fWdNiw0Uxwg13HM
yaKqUcO9NcC1VU6xCP166/bsRjcN5u/2YdT9bh0yWFpjrc1RaI8mM5p8OJTqaRcy
iEeAGJFWl/wrCxiyKLrFgNuVQs06isygnT14UIKpNIStRW6QeTO6EhE1+ANcVCOU
rlU+8wwmHjaUM31lpJp4POLSVM9bJrPb2tmFCRfiAqsW4NxSEcPEZYhSouRAM2ga
7d3lZSQFMHT/ZzjGFj1hC3qOmimTNhGYHxvAxegLrknCdDYcqDv7uw7YFlZQ/pNK
ei0v2fN9HVuBJ8H6kiFcFJSeVnf2Sb2Zcov7xleUHswq119DEiExQy3hOXpxStbb
5ZeiE6QvKHh8MG3ddut7AIvNpvI2zK2wndMWIx6t+ZEfjT+IAYBeJEWn8ATYjhm7
SicNYXN2yh3PtqwTs/StiLJ+IWDOPyLV6RXeRecDnoAGNWY7z3vOzlp4RX9+4f4T
Ntk3l41fcE/H2wAiGIIOKf0ts+9ncEElIEgtjGY7AX4YvsmGsYGfkoBrmREsXy4D
ldpSTZ2gyzro/50PUydckc7wSPeBKs3vm5lhlHiRIxP08vPzrYZ8e6evpKN8pq3h
FcBBtfdT46cMQy4xDKk9xVulX0C1YL52et2ugna8P2jYi03Yq+vwPkEHm9TavaAu
6LWIlNWCbQ720Tf5uscbFFgcU1F9zqOsc20KSJ+wlfLJ4geMb8ujOQhsZMg22ynG
skaFx7BUDLDn7oXgBBMhdntXTBNEGyCiQ1mS8NHGk+Qn7BONQ4xBHIHoK2UIZZdK
4C6tvQ/btGmpI+lX53RPHVPrTcjOzARXE3jp/1+42ZHBswqtvCnzIWDX/KNBt4m1
nHgb7p0SF3eOAAfzA55KJ7VbzHYJIXs5D6N2LU/vxjS493B2fA+s9Ejk5ikKcq92
gJcNYxh2eHoWLND06SUe57OE0VgyoT0ePXTh74/qjqikX6J7K8cCldY2zp4/vnJd
DVLSvRv1yafEKmXeOlSt05dXq9uA4sG5dJOvOuTTzYDyU84szxu83GE8a+cGvfAF
4l8JnxilC5D0ft0CsfASnTEOh+7YpHtS/r54fCegJrh7AG1VqFUeigIZ9+Hh7a6O
cIuek3aS2XeWzmVdziWnn4fgGfNeVJHuXBvR25kR/ppylbm8dY6kmcCBhzBI/vvz
7sjcL698heabGh7Jwh4phzQmC5CyK/QSDJMZODQ33ugIQp5VnwscBok9b0qC0PTa
yUlwuCS4v56smjaOQaIiwL7jjQR0Hb153zgZ1ydfvaYsz7aTvdWzZPPA/Om6HtZ1
w/hSRJM/XliQe1yFF7at9He3ah8SH0JBEAGDxMllt1bocRbrGpcsh+V/0JnTPMtJ
0zYvrEj49NaQAY1HK2+MjixTUa4LOjeqU3lK49TeK5x27Jr0Vfu0eTZb8kY4HQug
8L0g9g26oIGISWd9scQJ7DlR7yZ9LfeupdzSRe4yujKgJw1ukbW73MhoUbZ21X2+
1fDnt1nYIDUs+yQ2IubcHoaOxhYdq2dNg2kMEijXupcBjFrmjH6D3vz0KrbRtef2
Mk2L/EJXRQJFcuYCQuDN4rQwoQdNFerLDzl6Ci0PK6NWwHrRJTuC8uhMd4H7wQoO
tYWqBIFZfT+qUK2tII0WKW9wHdiTDb9/9eqBqUBaRfbeKRf02fWT1GEobjq5dN0I
sDh3Ms8yf/vKT2BmjSGDPYzty+LrdnzDlkxYY7n+233R90V6lkd9YwXaumDF/yfO
hsna2F2wciOLcC71Ulgokli0gaYzLHLvqRadQv8+DqtmZIixnVHnTZk1G4zsxWwG
HN7aL6ZAuipqTv+QUenTGPt7T2XSvBiH7LzL2Dx1tDk8ozTmyBbdFh6Ddg4ftfiK
NZ0cTxbNaQcCDUn/yXKJv3HUBXmlE4EkFhHThh0xSeabUkU61Gl1jDNE+HnCv8Fg
ILn8fG6bt42aLzZJwOGVx6RZwkr9k0HYJV6O81b8Z2RqlEh61orPRVysCHw1JCZn
MiD/o4Cvhy7EXh+HpSQO4Z82LPzpF+wCIle8CkrK5mJBTuWTNrl4krhJRXcs82S4
gGdJZJYGnciZbCOGG4SYwSQmh6u5PWAz6i9SE9gW4Q4TGeIIG2VanzDZw92IoYYN
GWNb9vs0lzqXqhVq7kSO6ex5SoPeyVI2Y2bQGc088fMfMEKED7nXU3EJyN9t7ZzY
wm+fFGMPP/CPDRm4tFOaRrMUpIuUrLqWI01mS4KX01qVycDyiHjQmCMQPOeFFqUs
UUGIE5xZTdV36FXhL4v0w7r2lglv+A3F+v+goNoyUPedMTlmBerbHDvIO3502pvV
oYyqvusIboYNdBYoAX8/ypUk8tYNw8ALkiJ/7dYRkhA+yqblQjQBwhiT5UMq7KUi
OhqX/P2ZAtNwSthiauzaFXfbxqK/GoqPefHRBRJCgBIsaRf3hYkxLHZr2REVs0tv
F/OBcs5PGnrngkqpuC7gnvdWxS+rl8VP+eKotupkXRYScaSTOtKv8IkigQLswwqm
tlLDo52Ht5JEo0E3ZhUFpicQB5qS7aQGAJrhKfbKjSy3qX9KAJejGF6bRxFYG2r3
FD2NZwyZRkwiZsFbLUNPkA86dK4KcZimxvqVZNvWCAKuQ0jmZ/COTmSG4xZmOuq0
jWabjqLcLPSIUYEQ8gHpSX1x92oSGa0OzQ2KkljbGMkP5IyNipje8jWPTLgCCF/F
2bIV0XeeMyVz51aQwvBX8sNevqXhh8y+TxjB7APtcl9uEUFDGldvGOqgVsnJ1Y4D
3Hj7gwxpHYrG1+0jYvZMMCjIkfo//Y6orkOz62ug7olmestP1XAJviW4M3AxIOr5
pp/oUVguDekBYQmHx4gzjGFthhnLt2V69+HW/HsyVD8y4UnBWXsmp6dhYYIMFfSZ
jZx38IKdS+Sba4BNhAyJ/tFjfDx7fOvI5NcoNVZci6H7RN0eWaONtzlRzLlThIwN
RqWdmowVK7fSnnaTa8iUFlx3EbOmCarcplExofYFnTtjVzo5aDWueCi/TR1rvg4Z
85gCvDzbsL3WYlmBtWH+1AsVKOVC3WHzNv9awcyXbQh3bsO5sQL4DMTpFoFGNlex
yfGhtzlopn5mDsusnS3lHHJgQrViKx16zxDMhjK5P/8P028x9e/rGzY7Apo+aG0k
xtIaNWTm2lwsns1eIObQJOSZ4xIQ/7di9YXuDjtPHF/zTB3XuI/UUzdZIPmswcOT
PgDESAQeMJJ8KS4JdtQ21ndJlqJE0RTbbRi7q3gle02bZW1ro8YTUu9xShC4PGlP
AJryw5oHE+eAkINQaZoOnXTpZCiERBEr/RdfTiWeZmX2pkj9B1QY/B+T8DOxU4Pz
86o/Hkffh8+h+XCtCKmm3YMZU6Aeksoq36rRWtM7KFagEayq2KiKw2/M2KQ5ydjc
DtJxueOpB6PvXc8c7+md9e/kXs8ZEs3OtGVgDdlPxnU68X4rGdqyUWGmsC35zpiK
oWiDdSQHw436fNSPtJQH2IgmA7E/BABV7jwfLCmET25XTFZtAUJJ2CCv6+yAJQ0q
eE7zo/QAIVr73ojGa7VJ8PAYYQWtwBhVmdx7ksAsCqtGG49XEhk60sO46d4loH4q
ULFm8LnTfbZVkuf6AZFKRbR0DBfdWNXyOEurKknpRgXsbfjqsmBNJZhsu8Nert1S
TMoOfMF8BfbcOvECESKz36VuM9e0fiOVrUnyqLOCtWym71/3W5gNX6hQPRSOo0/m
I59G+Sf+v/sT1r0wRoP5T5iGTURbRWlT3pRLkiKn2HpPzj6qOcOzJth4nxIh8XAK
gGHQJEXKWdo9NH5kPWQTKp6sKZ91wj5gdlc/kx2EFtqf3pyqWxMouPHLPY+UMeRG
Nwvp9gWO7Fo/++ViKUnNr8R1oQ4VOnHU3t9zNSMbSYrBCwCKO+TBmE7xzeJFhkaX
/TT3XfcSVqEG/Lpkm26n0WDIGH3W5RCEcHCVkhREFImGDGVehYpl7e89zWEjz6tA
wEB0VbT/HCYLvJIQjk0b17hOlyth8qAy6wy9c5oqSkG6KuC30HMDgGIDZrr4+2B/
6edMqVv2sOLfIuhHNXTBc8rTEn8c0cExx9VCPZ77UzsLbvi6VD5Zr6g+AAEnGOVP
W2tPAb3evbGCgv/gHWsrJzEvpIP3obJbZazPMe6zI39Lq50I30L6o2ZaWOeAsunh
oZh3kkXGq7ytU+8pIbtZZxqnfonwypcXGw072s4KDLedqQkjjD1+0LaSG5MpvSu1
+00vTr8fNcIxyBnVCY1N84HYxckFuCsJZsUUccDeEX2K/wzy7/MvBTschRQ4/Eov
41IXt/lZaYgxDrwGsWGWS1Q3j3j4ZGVjAXyC5GVFxHa8INSDLi89z8Bg/dYP2php
yUIuBJiWMrmksd/ROOd/8BC2zAyM/Z4wFLAl/814KSvaSPjuQY8tP52nCDRTS5bO
3fVVRb0bRkOfpvzwzj1zjny6FWOqTYqRGx2Dit8J1KTY3wPktW+ZrQa+4POi4RME
I9pAT8u7YiFP1hMAn+vgaomdojadm4eEU/yDNeQUp8o3/n0H0OrFceTPawNas+N2
6K68kWPy1+zU3gFLnffa2AC3MCikiJWaxBi683ggaoQljK4oJct5Bev/bxXy7OMv
FGo73GLznvl9N5z9gVUSeZH8SMzOgd6MxtYzSZJbu3+SoNNU+noXcXw8n5vSy4pc
xOMYoUsiZn6e+dGegOkC2YDxH9RfjFEaZ7G0YPkqivDb/jFBG1m1kBzCtMJiWs0a
iyVeCBGePiWEcw5hHm12FaC/ChJdOLLfteBFvrSZbzQUTPlv698bMXCuzVRFUQkL
qhH0VTAHC1naqC9wBIoFsYRSXd/T8fZZGnHIBOZej5t0WPNDGobgaa0SKqShHISO
P2pGOdVZdmj+FFEmcT8hcCGvkmtA4pk5DdU3Jp3A9M3ezjwwEFJMfOVFH7VKUUk5
rRKe/csVh57pzzXLqDCDMY3btqzEp7zqUXdurmRZ/NJFaUFI9p9CF09XXt+11/+U
XCzBlsF2dJM+GVdMHtCI9jmt1Bh5W+rhl6W23/2hU5Wu5ZxZr5H3sstlLj9UK1Lf
5XfbQDv8vzxXv7eDLLoVyzUslPl8rvmE5FZZWvk9rIgRghXboq9YmfH0CsqPlpoy
ZLA+EFZ4cXnMfGXNpjjACaUcxrAmzUEmU7vaUv3cq+S6D8mHRvsbez09wLyBK/6H
udzg6MFkdvompdX9Vj5l2QChm1Ce/UBw1WvyV4c8nbGgOZ+SWj4gUE/UML80XuLq
PYnZOpBxdheudp7lVPM4elzewjiTDAiah1FKjZVmEh4KriK66UBOhCz68jjO7cJa
Ng3NUwKPqdEOZ5XzkmK2lDRIp1EEHHUH2zb8fSeSt+XHHha7yNXUmeevIA45gQ9W
uLlHIIcphZ4vEJveXcb1aDI6CuTbaTRZ3NLgw/FgWgJRSpwpza9wBJ76i7phu4v7
QAByrpsRmsMiNLdgLFcm4RixouTE6Z5hbzNlhuUNPJ3VgqmuqZf94QSsDNJlfDRb
tm4ABD+Lvy4H+zzINvKrShS+RtWP3z+NESagtNm9Px3xMywcjzPZD0NNrM95eIAK
OGInzyENVSU5FPVIfJOZeHw7K9zz+zSAmdzak1FHNdL3+8JA0ZA7mh+kkS6mlXnv
8Hhcp3+ptuhPCMxW73WAv+eBvQiXaInS2qGKW+XPZk5qMYEqj0ZF42xqX6BDtE4O
Kc1yJfqoJuatjpIwKo5WMxxb4wrCIYJu/btO9l17Dpqmz1xItb4H6LdVbZbmYhcR
9jiW4iQFRIznRGg/z8sLkMJAllrMfKBmkKVqjXC+gYI4El/6PPqiKdVYQUdfAgc8
QLDycSQ/BrGBTVLKbQ0ca0OK7mOZhmSKr+B2XFdG3WXGFNsra4g5irre6PihsF62
Ibd18S/Vyt1J1Cmk6wfto2o51KDGoMbc48JjxFguqHNRidq8uy4nV8wfxDaiTi2k
zkcZ9r68XkELVxT6x8GIKXsajbf9hyq69Gf4Jn1z9sZVIGaRRrvAgqNyr4oj9Uv+
cfeVH6x2gmEFejM6ph3CXu/BT2vPJK8VArLD4SuesuyFrlo20S2vS5DR1v5qJCak
zgdA07xOYwDUu9sTrLsgpf4LhanUzf9LibQG078+3I0Qk++/0VtbDySpks3Oe9Nj
EGsQh8W84TqS7eaJH363gFt0WB7mQCWFPN2hT3Q1nkW4bZSBqPrTuKzrDdb40pqh
Al8zGptEv8qjMVAMgajRcwKOaileqxHNCv2Xy3wEGRm/vlXuEO8L3LZ8QTPXhG/k
Wh5mMzzZ2j2ceoMFtuNBPH9qPf+ATFKjnmnA/x6sz9NaqJ7HbvpM8I56nR6ODX3M
Z8AKxvP7WPkzPrTygPW3pthUWpLHa2xidZ86Jj/O21w92QpmkgqfUprbkSoEKbNA
ldg4J6x68ANQmQvxALmkLt0VWFrkiKh2po/STNF4ODJx5o91k85JI8E4/S/Z4eRk
X9jCxThXscKYFOJKEJUFWuyO2qQGq4kTdF+bl2DyaxG8Mxfhc9oQjzdVP3PVkfUN
sNZ9w2QmPvQzNlhGNp8QQVLokhw11fjJuXORTJM1jOfMCN5HAWHJCpCUVK8H/hmW
ZBn+CpPtlHNkIJHPCRfetJ89A2FkvRBuGbcp/dsXMWzcmw8d0xeSKA7AKwmuOJII
BnMpFmgWxxSn0XWCQcyb/5G4/6UJswQqsBEAy/Z5oTA5/4TQK/lxqGKWQi51h0Dn
Y2cpzxy3l5pSMTHi7R4oUWENPW1HVk5SQBi0cSpQuRaP4uz3qMXTTajPA4lL2lEe
k8dIIJbXb1kiejauVmL3w9Q/rxOg+6iezmpC6hz20RODE+c4SOJ9lVJSsORN6uxx
UxgmU9AmIuZY5M+at4zUt696U1+vZL/vu3ZJujHUZ/NiS1z1005dqHlLwVgi5Pf/
TpJx2wgov389Tc71VX6BBls+Ht4xjVgXBCWmKJCMXBd+nDzve+ub3FA9jarxz01D
Kmg6dJRigddxeTHUjGrmwW9wZoC+HKxWjHuRU5vkGJ593Oih3WfYFdilJb388tyq
6GUwLPYyiTMN1NDcHpkFcBJppMIKUMRDs8MJpUz1NPNl0+aL6eU65sAK3fwwytXR
/u49P0BsWf0hN2fLSk92zSYXeXhCTbRie1rMoMcMF/n/hg7gfiCDcjPP2+3Fu7AL
A7EQT1vjRSsXFCf/lCxJNcurYjAMatKPM6afLXAaSoPXbFkC9MIU89HizalTljft
/8uCpiUnfPA7cIvFSIc1BsANJ+Fzt72AAnkv7hCUrytH+gCSS9wE6nEIMj3a7zit
0b41YVYLM2vaTs9bolb1QWczXpnfM4S0Ppn7eS9bw25Noe+ZFXd3fdwNRKvOdiqy
h91q3OAbPhvE0042zZ1osq8QKWi0T2JCX36RDyd7nBeTCFml71xE/Dv9PFQ1YAcO
Mqr973he3JPr545e5LLGvEdiKGyFVT0+cJBr6pw1o+f4s9P42VxgIukjRyxL6E0K
bjdKG2SrJp79BDoYi6kcMaja7UYTudeC+UoLVjmZob3g+JDa0AKBfA5i53vSbcsP
N1GhiYhcihetbSDcRWClQXzptNEZBOKcaM0DpLkkiQtsnZQdfEfsHM2lV8WumIEl
sjJYnv88SO5IZuOfmgQQkAwxy3HV0xVj+FYtsjhzPvXEUdKyna0LJHTKdQXXloMi
Ws+rUZiNhKShLttOnF7opXMzyp1AY1xzG4iGiSh7wadWLzBuS+vpn4ErmWauiWLl
tVXIn9qYkbzObcXQaYKeoG9+06oa3uDaoNZbkLJKNe+8GMaQFtj9f+4XQw+pF2Sz
MTqI7TVa7y5N4pHDYlCZL9p9Bq6VqhoGLCK2YxMyUo6Z6y1X4Ypkbl4rfQikjpMO
HnjhJ+7eIx5rU7o/A/TIXyTOf2F34qljeLVIbI2zA1xtFC058iMWuF0UeMNGEWWB
yUbZOWkrOKn7dF8WrbmOtsEphqS8tFX6uSQbxp/YFEpky+ge0l8FYZDA7cUxkGQC
eL4Fx/q8zdgZwHtVMtR0NB6mrfwXeDguYt1YxWsFOgmkvkiSQvlAls17zrD/zBq2
7AR8gA4MFV7DFD2YjFSt1kwjmbTy+3YtgNUlCv1JEXL6JasJEvKL/YvTjibcVdVr
8NjYczVhu/KaKrTY4vSS1vhngUnS2yRLwJXdxBtmCupjmwoxF6d4Ypr29xhNFUGP
3iRgjKqB20aOVLCjSVWAngkZsKuWCRsX6t64+05i9GVjLRhGaxtWjw7rqLljrQsW
ey/6ZWHkRXWyI0g/7PXKSFm0wN8xr4SZw0oyx4erz+Lx0P+8t1acxPsa9TTCUD2P
DC7kkCPXn6BdzeITsiUBesjIyRxHvUJpDjQU5TNoEZ0T9dYV38Bvj2xiCzNsXLAH
FjTCxETMVYi4vbTI0TVBWPhYF7Rj2eCgpgvSVNWgWYcmFC2LaIQxmrfEcg144wXK
LP6BCblIDlU7sB0i2zX8y/8hOGrygajUy3XKZs/QLJiMXv4XvF1YsOYXBZuUSyCl
L2JPEEsv9+8kO4MBdpU9ivwtV1OuRW6bc9SxeBcsd68XQa9oWqhBl0vsUWz3gxIz
tKysiDXOA3aU544WJbBuWjGCBLzDjaAbh7FaRDQh14Z3lgxxKrwvt0pOYzayHjCr
Ww16CE+FqsTG5SDEhJKTSUc2pFw1E8c6W2He6Ju/WkxhbOpAVXyf6vcP4a/MRO+3
1GaFCYZNiE1XzDeioZMQWThRAjb8rMrtjXkVI9ZJpwYFxSMgSGl/oJRfKS3POZpJ
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bnBmVcce36ru7ZaWi31BEkrTJBolpwIyOYHdIHwVfYmd8YLy4qCU6c9511PuAjkF
ETZEB8m1JmzSBxrfbyELsDhyVbr0bah+owWBcB/vYgBH5Rzefo789hu+Odz1XsBT
vQTm0eEvg+qHAIpkPANIzJmNbdNQaiRU9lGtdD74yXFkLDzUmDfOH7hnPPOWIlD5
1We4W9z2x2c1SIUUvxz6PlMv0Ye2YQwkAQ3gbQIM4tqd3gt3zA88jzwRo1VFgRXM
58osrUL2X1AiS2ZXUi6BdBxX5SlISMx0l9a19RNOs+ivMvfGGn35G9VhPYLcDA2p
yJw8uVE45E9gnMAoBel1jw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5312 )
`pragma protect data_block
e0pABY1+DX2DMB6CdybAqDFYuqdGbMGCNZgJ5nxP/LUw0fCTABiMKyiqveeUc/ia
kXdQ3qXI+zrIMW+EHREQrcMEDeeljDV3qDjNUhqcm212AH3xMBc1c61r343VEAUl
ppjlkYq08dXPt6wrpfI1Hdkp1cjbo7ZEV0+ykU4f9ags+KsJ0AezObk0JG+VFaHK
8D/Jn5JipNyb3+wLiRT3LeZ2xg9CWL6brit6B0Z9xJ7trLG6STYVF2VvMAyUYv5i
CNpxy3aVpY+VFCISSsvmOCiTuDPLPIatAc9X/EvjmS7v8GU9b/7G2MOyROjhfQ+H
IWPfQRltyT1vZDvsVBMeWXdQ+fHFAekP5CFZs+FHtZOpROcdr+cYoFNtQFFBlsnW
vGPwvD9u2rIXSakLCL14dFsZp6k/8OyNu/MjkgrBISRcQsnrIGqt74Zvoieeunty
/ULbytAz/N2dr45yghRo4nE50C2CwNn+xLTr3c7zJdOhwLiIvfy9jK5SuOGFcCiu
eca3PXAz0304Iuc9hDB1HEPkf4gle/p/fOMLm/fsZB22Lu1khbp58avpvHjeyCLu
KCXevX1u3fe8ItTB3K4htVraB+W+nBAFA+qCOu1mLLZUUDuVgGflFQOGjQaoJJYD
0uEm+Obo/XTCVvb7qx3fsDFYqjGYg75A7D4RZGGof+EbzT0ctge2sjCR7TCHN8Td
xpBOQ5SLCn7KGDtG+ETAHUgV9QvvJ3pmtHg1DhDUD9o06fCcyfVLFyT/Ym9htqOw
QV/tZlV6LHJlGQVz0r1rY/wddUwiv6jK9d85bF5v0EI1pYYwioXpS8byhyvz8DHy
s1tv83uEUcJh0YE6eQ+8VB/MaONXTr110u0TvUk4EhEMP1azfS8k6p6eaeBSqEtc
fX8TdqB49T8w2dxDzeWeIovnne+AIlwp4KBtDM4Fe7jFItJqHAACjSkvWCpu9qou
uhV4Waw/BZ2bvKzklGUBonPtCh9nlhUsVTVhCKDZw0JQ+W4a9tHqQwD+fEW+DeR3
v9lDKxZ7fx4NKdTFtJn1bkDRo8rzsdicnKUSQqsSmPuch6WZpdboCloLXjlrMNcH
vQZ10INcJ0brcXgdpZdNerT85W9dKH71xKptGhazKNbS38q4KFTcYW8HFyTg0vJg
pHMQ3iAM70KTlMFDIJBGuZN8w4W64qR64s/rSAV4pIjBvof+cL5/9V/+XHc0yZRH
kCW/8vNM3x5lDz9eIhlfAknlPN/fPoApv6Al2hxoIXTW/sa+UHZpuob5OgIojy0/
Pyr1D693hJBjzmEUSc/6Flq2S4E5CFRTZtrvFUnAkm41obYhcJth1B+s2x3QQAes
uUGqt2f+agiQfY/Ucj5qtpzWAX3tSdSVypuAY6X7LUZO5BE/9xxJyS6fyQMUJiPx
EFYHxLiufcFPF9zBZmgXkkN93vIKQdY3U9C19aQ94hR6uXi1o4oHNbvPLha6XJ9t
HC9zooB+nquTZKOzn0sBgl+A/RtMw3vdhbpJnWtmWiQISOWg6CenCHGsdoTJku+0
QHOEIW8/xYWq+y8og/pQS98gCye4h0CDZGzjNq/vtBoYYImIW4ZK+ws/IytkGO52
seWfExqUQJL6eDQI+7q/U/cVI+1IZaiZIp93ZyITF9SnY3AWQmZqHo8wLPvAqazl
7GHVKSt3uhk90N9KmnzEf+XOBkrOAFfcsvAbHOZjHbav0jzxaAw8K+XwnvpxNzsv
FAg393mz8zyj5Zjkf9d1Zyae8l6PY9UllwG05OOJFJq1cn//UFLEVnPVf8GGIWPI
AEHok3/HPZo2m7RUrg71wbAQ7V7V8Si8TbIXJ/G2vhyS8wtdPFbD//wcbeo2323E
WLtIRgFkC+hfxX7z717STbMai4vLLq3AJHQx7uoyVax8GRt3UoRCskdOkkBaIHKH
g2Z64Ibd5/ggubNW5HgNTpLbyqmkA7o3PBNOmyajMRug8qcMiWNfFq0crw1ZVqw3
KRdUgOrYwzdrK6fN+FTKG/9XTdScmHAA3JrG8er+j39UxW6O4x/Sxt2PaUQhMzKv
gYW/HORxLlcpi6vslWXi4yym1RHCfZQ/2JYTphktyR0QEnRLp6dc+Ef0B3FxVCVs
BmrVC2SvCRMuSVWYzT7rBsgJ0032sVGUYHkeCXpcMeMO5zOplFoIwuYrFB1PhVOs
o6polHeTPtQHO1tyWXIWbDmiEELd/KbiVsFiKrW49Smsyk9YljBxN8CprIoGjz4x
lGJKOvtP35dIyj7CKAcoA0MA+ZRuAr4jM2wvRfRveHwUS3uwJEOBRztSp/hZP6fs
58UZKYsTtLWonaEidnn2pfsssLFjapjf5md5/edoKNUxn+eSj+RiaVnCWWsT0rJV
rWasIMLQ5MUlSFu/sgzULFe9wg+4WLSQkPE+44eXkAVzUpAFA/M5Y172avvZ3aiw
inWq30Re8VMyohFDSQ+TLnquJItjPiYai10cs2QvdFA+TsDKMljgoSHGu4GZv2a2
I9+4oyPDNFLPzsH7eDZGkaAUTagBYWvrFI2KrmemVALbtb323hkapyxrffoO2kIo
oBfjicNCYmxqBZWop0QIhXH/ep0jjN43F4twM941lKPtHLvRShWRMByQS/A2B6p4
1kgsalFBlW3ZwivjqDWrDM6vucMLeb6SX26DpNfsgLYMwNcsYbS031ZxYGWr9+RM
JCFNCTI7sjtR7XJYZ5xw2d4UeASHmwTLAc2CRQagMyBKDbyVissMoWcOW47ZCMay
lM3DcqOhbiaQhf9+H952yEoci66mI4HZs9/PKkEAX0XdueQEWjBPQCrdxOKxjAlS
SYxXj0+rtzDUYGs8/4eAXJhDW3rXN00nv8uRbP9pPKMFg6hNSv0kLbpZP7nlZ125
cKgaxhCKOVozC8D5EWnkP9o4BVK9V4D5foBfaL7SptemTzozpbL/4475X4fU30pi
pag215RDKoJq4Y9s/AYXon9+Qm6Unbgpigga7PKSGGK2OMieqnjxhI63bBtLgmOs
00YWZ1rWElS6Y/YiYUoPRk1w3kv3384edvIs08JVvWoiLe/A1vVpL5f31Qrzzs9l
zhu+BpMl8UQWitF2rRGTCwjo2cmyW2LyzrzuNPGW2AOlanyG76zx89kDP4qLn/Iz
YIX3wruRuwza4TE6WRoIP7bBEO7rZxZmUTCpYJzGQ+joi1QmJdBi1vmKH6SktbUd
zWoYe/ZstJccW6cCLmrw9hH4m03eI91+PbxW1QM+5fjbqRp00rdH+vspxD6iilVB
SH3ZiVRzmFh5DinLU0WFU4Crw7ccy71m+4COAR/Nomb61+m2v+hd6Ldx/DlIVYFl
6XuTEaZBmUmOXIRrNyU+c3MMhPj7cJOSRHbtWTYZEgeM0giier4ngfQsTBBkyrKx
FP/uNXog4MXjymep/r+uyxneLeAzXjcNA6dI8TGIaTBr4CcNTMuI6n4xdVXsTSA6
NZKD1vRvtoa+ld0m6B07erbys8E8hzZ1psK2foA8mt6y+Ta8CMuDppsUE05ykTJu
cKmPEmrw8YFnMGUapoNd4nG10JBf7li+CS2AYKNajAYv0ho6TD8JTHVjdkHk7bwS
+WzRyy0lSeOk7F1VHNSIH2U74G3fVTJK+mewsx5fytGZEoYyHtOWqpYiIDRQPMX4
U7gdTjZLgsHXslVE4qIMFd+Jmrpb9p4gcLgRr+eBhULALIB6VY0z+cJvmoCWli8d
lMULaZ6T3RN2EoiyLMU+S7D4AsQZrS9cyAdzmUpHA/JAZHYoJBnVlvrXaT1Y4iHs
Rzs+OHQdutEbVZPPIzfHB89kHA2ceCmYW3kiyLs0grYCIyk/U+Obk7PPP8mxuxxP
ZZVsvN1orFPIXQmmPaoOE//E8nPT6MEAWtglgdTa6vOmRhOkiIPoI10p4opEK90R
7YkZjiwa+2N5jjpcBqkP3/sxPURmo4no3JLfscP3iIh3Bbk72o5tAYi4OhUqCAcx
FyJ1GX6j/N/dwNP40X96FypyGpYy8gMDsWRtnqcYZtOOACxDmhBUVYvGlP3LO6MN
klN3XHCZULOmnFdmxOH+VbcZlHWF45AKqmJvr0WQQsRPST2umU3iM2AZJVYikojI
V90rijv3mMqaSdBQZeAp7wnTef0USRm7E3pII0mCgj4ejhhhlgo6Po8ye9NZp/li
LUwmC1VZ0bmvk53okXPlnQxraztBNdnus8l7GJQU2IOKIA0mxAZ6MtwRuY8OZ5A9
wbvObEEusZIueDmzCDuu9VfoQhVOe7D2qqhHOulSvE/dnRn9pC5xprdnK5j7xxjX
T21GOunVXvuahEh4w0mu2C0tqL04Y+ytVD6O4kgGQrCmzfo5vWxB54taaWEpgBft
+Z7c3xCWaHLQ+N8Mwj5sl11RBA8iN8b14b2GOFDBLhRfQGZE0xe6H+2Z89UMXKPM
UDQYXu3/E+Cth5mmeQzPPBKogUuGplzvJKwHO90PHCZrf7osKtzc/b+34QReMls8
10KHT5TFw5C+FCChy3xV2fXreoZfPpASXSwIJCHHxTGfJhPJ8N4uk78q6O/HgIPf
m3Q0RyqGVrajl09SIxoWOPs+VUNys2krHwC0xtbcQBHf4qVGzL4LXmEPSI8d76MG
NJoqlfhNsdfE4f0Utjb1sKH3ERgPJ2eJezPT6xbwoBY2new8YsbDBoSegALWUKHY
v+4BM26jOqIZpLUxsZkNQVFu0dKLDmgisPaOM+L6XLJtkuMZiMr3QxUT1NXdPHne
8KsviKE2ugGZRYiV3Ey7b2KxA0535ZSVRc37S/Xyg4tsO4IaG+0dkpmwHuDlozua
t2rFJEzPbG2B/3mKEizdCFPppkFzBfF4/f0uz8vxM5jIPk9nW3Cbl4LDoKqWR/+r
jo3vEIIiP5s3vFHQp2xTfKMr/4GOLevrPIEC7YUQMuzGuV/ns80RAqoLASS4Hhd6
2KkovUjFlA/VocjhJXZh+HvWHoMEP8sz4H/+j6Nz7B+5VG1DAxJ1gjZMU4G4OGAp
VD5YQGpiVKPz5bb/C0pU3pjM7jP7FJj8+hC5RP8gtW+0xr2J3uYFS6Tnw80Vcsop
6gkZ9knTl281iXqwMbI+0iYVERb2PakUMJDobQoR5B9SOJPOiOehPRPGWWpRVirZ
cC/sInvsphdoxcIWlMEZkgh36+nMXdD10RlJH0DCxJhEQcAVPrqwLPVXjjDH0OSJ
srdZWpSu8Gn4eWp72TVTPpUpXvl2s73RDepIeiMygArgQrQvFdlQuM4lp1Q336SO
QTnYcYxXH2yJBGeRCTGVBjwTkaHwIwsT6wTYG0qdU1/fUuMnaZ3TtViGdRoG2FKk
zUXrcttrzEsSyxRvplOzifMyFh8ZTpEThAvuYs8LAsfFGgdiHGEul/OeKa/ruhj3
Loq1vsrVMIrhI2nzH5bdTVuBCwVdrPTgYjhnBWFTunia+LD+er4Bbu5Vnuy8P0pm
60P/hfBID34x7s8JS1xgMlRf8HNOPJCwKJlxSiE3Ln3LBSKBGonwMX6YtOIQto9W
3SO901QDnv7OnYy7mhlp6jPq3h50ze465ueI7bhXMjZ93ShTzRrqr5tmSDHQu3NC
08Lk/la1ihfEx7YyXRkTvwpRC22GDgoxGSWXSF0kfnU5sAL+are4SO9/W24RQWiA
7KgMwDGbmdMnHOhfYzpMqqYxL9sRnWfZeNHMaSH8+Y33uIr2KgPKNJPgj1Q879QJ
Obu9XNFsNXhDFAR72eHG7/LseCSiadgRjc2PQaTQLyK2tuwzFvUJ/+nyUdOha7Bp
9uW8wmly0EV1XVIEmKs694EFizX2yxjTRO4kQN/G1U2DS3haN8LUlO0sQC0/HbxB
Dx5bWj574yu9xWsuKEMffwEo/FhGNNE37Mb+CiNhYnARUN3gEreJWv7xYck2U1xq
GvvxUwHyJ3syjroQgAa7LDB2GTpb4IplgSbumQDRVoKwgh7san66ZvMj+ERTIkIR
f2/I0J5PgTjbGy3njmzLB5KgiceZXAomlvbKMugyXfWXlxyNeanFKdifLNlTkDtj
zzfVwLOVF7LVwd2ZGxzM7N4XcMJkuAYlo775mGoHOyW/826BiW52ocSULwD1SpgI
O8JOtp555scVJ6RRpSMRSr5RKRGdCgVhOBFZpwFLjcgfnfL8rKRa9QoQkn+3z/2u
YQVnI11y4EFfH0AzVtbok64G/MHRlcnB08QgY+KNQNMVujWgJn9E5uuT7w8K+FzD
27+3FJ7d7UTOS3tn6GdRiqr2Ly4wGV7YST73Ly3A9Uj+wV23mBkQ8sYnrEk+l6Ww
4LLFnu3ydWAuIUODHowoL2i+clcI/ugKA9swN5V8dh4L8Rl8rqDCHR67Ky44bZP0
4MsqVA+KwKIfvnclwU7QYpLkyx+EfuT1/XAcONGwe9H2/xlMkdZT0WyiM4CM1W7l
26lhc1W03kt/h6D8RThXtgSaK0GHlTybJcxIRamIYZBmlsinGpCrC9uAD8TS/16o
hSGKOAJ0BxRxmNhi2pO9ojCQPj2ljzX1Tlt9iE6CN9gHotMt803DF/eUelcWFrsy
Slu8Xr+CGVTIn69+/cI6iOd6P2uD1DLDh9jLmG/+xcqWMbB/UYrVimYYSOKbfSdw
fHEYCa0Joyk3qEhpp0TGdOVVmlWS5leUuF2XLeNnniFECVZepX7cicR/MslUPGzz
D5Rkb+zOkGDeDSJa4mKLAFhfNmwL/mLjN4YNbF1D+RbA6uybLRcdKbdfIKkC7SOU
J980JN502rjbj0Vs068lm/wxEJP9VBvHs81RO7DFIl8oWFWGLwluy+4m2n4Sqv3T
yMp7UnnvypADQNVqgRlHjZXzQdaURKeQ9EqGj/c1JJsYIQdG1dFwFaKjCjVms+pb
8AtkxK5x2lkBQMRoyC99woyyDQOHOh4SFCr9A1IvO9O0LLzfOGMQIPCDo3FcapaQ
3T4CWaflQ/U0B23RL4Fl71VaKrJNfVnAxo6gEaAsKzfutWO2whYaOcQ2lgm7ztH1
slVnRjy0AFEe1zzXm8b4BT214NV5RjYxdDjJKz2QGLEMYGT0nMzXf1lJUhHsFFie
j3W8BNMBxlSmcCePu7IqwCtiZ4xEtGIrVgRbCqwUOKo=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
hWBSR14j8jG7F2MTw4h2MwcBDEVJASKbCt7MYh+pDPaa5+RDF9XQIGBXbVwYDnv3
mk64qQO9M1LLDXqbZO/vxb0gjova7dg5fWn/17gwc/D9xZJkjNRrT7NvwMnXWeyM
mClNx0WCAMxekgoZAxFLSjCLClPlMJa1uLjIO43xHgnpfKqgsP1ILQKWw84NfWT1
MPSOxX3/h3yLA4ZZTcLToT1/zJKQ7Tck2tXXyXSjNLw7Pt8SV4v05iQM0UXsDUKf
RE4dBLEl/kCVxDHp8cf7g63Xfl86A4vbovpEv/bt/1EkCclUWOHSZ8Usrx8VdxZQ
uFtytf4uNu2MgHITz8cEDg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8240 )
`pragma protect data_block
/Wwbqo+7SXW4Ou5Bg/MQ3nCu87SEbSLqyOApDEq/ZxueB2VYo91J1GcHigvznd44
PmR4E03XIX2N1gJOTzzfvqcH/q6d3mHlsDHRISlsNqPh5ocfUE0ikkl382GzgiX9
IJ1AsS9fAonXeTjzNCGxvvGTiGEXeAdGiTqFWX+z9JD0p1BfbQFTYl2jNqkSeSMU
O85x4f6jRS0j1vxRksB15L/lxt6PuDPj/M0w6Ui2gU+7k4kNy2w/YbewwkE6JPf7
3hoPfQFAmZwOp8NfyCOJ9GwgjsdCxqJa3viIV/4US4yBWFpQMhiSGwY3oUF5/jNu
u2BplevMwPTp+C++Ke2CJWunitewKCkaAWoe8qHpYbHe7s2A7s0UK8m1EEaF26h8
7BDY6mtvUzTVE7pW3p7uBoS7Qk6/kzmec7oHPtP7rnvBFs0NvLeTxhQEOr7SZ2ER
Agm3ODklH6UI18WHXc9+bDd6sJOUfnTUPUs6No+fJ1fdkKOoaQwNX2jZEEhWOWGU
xWQb8fpA/cmfde+nvLuPLsc3MBiJpaSF3JDaP3RvFHZKotKLiNk++6yLOgMHb0vv
u9Np4nfHZVjaMeZfz5Uug5JPPiOQW5ESkSa6RBQv44UJcnES0hZ7R32KBD6cTRQT
Rt/0lV0xLvVm3opBkECpJ2RmmH0y8nngNgPEJpgqMDb+Q+SPzFXBQ7UnJDpCCTMU
YYx2Ggi1Fk+3xdVbILVwPdHtKvGja3ekm6F9hTOOAU0DgaQp3e7ne6ruBHd4Fo71
KYKfUECu8bEdm1kQOFm7prNSQXgIbFunvqORm9xfH0r4TUOy6ItQKeb2Z2sp8AJM
Z5XlbVncFBVnleL7I4o+V7tPmu0pyQfJQBq2jeKUhzMAPzL4+xOLX3sIrShG4IYf
SK69DIGTF0jjU0XVFQf5tnffale1vQAXSXu/glmqDCZx2rd+OnVSAJD/RQLP3abo
pg6FnLmoFzI09hNAvu+4LyzFC5X1PG3ToqTfIQZv3PoHHSPf4mTJUB+K6ubGykNh
Ws3OSWKVE+q+cwjacVqb/10ZeAC1Bgzt0VHXKTFegbYXOWnVbQeg9Fsf0G5vsMyK
7/PlIBVH6tc3P9sAqvDlc4d92z4PH40Wg7HZtWcPYcD/gN5HYlLp783Wk9BwERDb
u+q9Wmcti5zG6ywLmPyJekm/XS9mU48hoX7hbwODa+smzvRDOdD/g133r887iR8K
/OKsnCa7t54zLthuCs2Pgxk6vT+Cx4mr7L8sBbe1JrBotlYxXXdc5kx8PAhRCCmf
ghRpQZ2DQN7TRakaYRWWsKNiA5aSxGyrXdT1MBNu4kn6xUxh6hvPgw4ZCsMxZiC6
N4O6rmleJRNH6UUT6bsFJBdobrVw3j2xGt+TDYsLxLRhM2yhv/4m+pL5glllHlb9
7O2iAIWkzwqKEt+gIgt05ZkfxQ0Qd7xNMmQv305o5xM3azf7nNyFOzJ3A6VLjPjs
4uhzg5+BJzv0GHvwOkjDlQfX+lMAGRY6ljTAkaMn6r8RIXx45OomH2B0b2EGGoyk
BdwehOWUQG8FNCI9BlkspdfjXdfGXXS9X1wyRBFlXToOsllLITheLEOFf1rskxoz
vhYYudT6yGBFfRMXsayM/EVRcdYBHXSACnv4ECzaaNvn3IYkf3ndx63cHALIRqBH
iazz8UeEUfUef20R+zYRV2DWbIDSD1/ONYhsy3BFJu7zUfuYhmz+vTdTbvH+Q+wW
Sa21ayYdAYdK59soFhvy9cRDo3GF5n9UUcO0Sa0TWTLEfVQuZ6Pq9iW3srIKwQLN
xuPSuNsd3HbzReIisiiNC4ZORE5hlY1oEzojwIidBiyb07E6JEZk/tLkS/6dXw1m
ghPvhwCJAhanbNjtabC1ilbjQ3dk3aZRPUma90so5DF+uOSYXS07JtvUqBjbsqD5
oXjnWyLERenToApMjupq11mHPlUB5KCHX4FAX/CX7FdTj1L2p+XjrNdx4dw7XKJb
4zQb+Dm0/xL5SapCoBKgyveQFf8ljRXv0MP9yoHj9QPVdXRv7JqFM4LsG3emTgIj
OL8u6fVLGa8s0CxIAvNH4E44ct+hb4d8eOfFrGA+FZvHyoO+VugTXwvdBY1M0heM
5X2jFCDgbWItmFW+yMPYAUYB80PkwgmAqsB+A5TqnRBMF+BXjjen4dtD37kZPBDB
83TpypGisr/1FvhEL5UhO+vdigPG2GiYt+wJqE7RtRHdYaYVFbguKx9P1milEItR
tJ/FhuivzHB25da9G13ZjRWQOecVFf2Z6bXPBwcLa7Au7rTftQO5JSa6tif48Vmg
fcThy0HfSyBC9fTVpyvUq+cN0u2WrIjB2DZMWc8/t0ijQccaodikORwCn+r7ky3F
M6EhGOG2SQdHzn2ai+uI8a3ndztmqKT5WKFQaGcSKeVQ+hDGt/8gx3FHJvNuAxpY
DaSmHgJ8/z6ylcMgRT0CIWeIWpquZ5J40cDnDPdDdMlcMo1seJ0KLg03zuLlBxTf
MNyr+5AHnqI2UbFkgx7WU46tpsBq8htqCIS9aEauvmPdtJ1ecY1lc0jtnTsYbq9y
MB4Uuff7JK1VRalLkfiuRXznN33CORpoAHk2eTiDiOl1YO6u1iJJxHUkoBIBYoTX
FA4vIJDr0X29pWJ4q+d9bBpqBdf61vnjqTLX+NgaPzretHpLz0SgAcoU/uuVRylq
I6LZucQmczlXRJbdkjkWM/klWUYXOHaai+r4be7vqWFThG32EC3RH+ZY9sJhdse6
cRSBNOFGJxyulJM1IPewmvDRAgbQzB7V2J6F0SXjnElvyjKkWt9fjY26cvMCgdW7
pvwnR4oN2PUKFQC6WBi+MrC6vjoH0pGeRNbMItzxpI9nzHMlGff/xHgWgbBrjDEW
t3ZxW5B9gSi8kJWun0yQVP++6hny9RKcLhOtNIsBzdCwkSjXC38l/1zNgeeYrFwb
cmdv30O1haRXdIzMd1vO4iqVtO+QsfSCFM7TKA89KmpUaR4v6EvqeKWK3VNrzLnv
Ik3GtuKpqFUMgK8T0lMI0KJhwnMDS3GCE7ueTIlO505UDNcB/4oQOBSntoz0mnHb
Ubv1y0s0iXyGdCXY14vaNzru3bXXS3JXOgrZamw6qKldnn8aoH36sWZKqKfxxF1M
OydTbtMgyWL+KW9gGBlneireKSfBLrf0ePwd6pfA4g4E/NnBz4Uoz1g3tMsGzBsa
+aebXPbp+JhRmXuvX2aX+sbIBxgmrgJWzYtS9zHEN8nu8inXslaFFgiEUhUiVAHI
JK4ajPMwxm9QXPDwGTUGcM9mkADQo2C3Cz1/Hv920S26u4Lf8YZ2VfmvXtGTtEL+
Nl5XqAewWsXkOyG7QBuuGFdv/ZO+89U7epIw3LLMRnpKYObuVQaJPGFeocvo0GUB
fUZyE8Y0YXdTiMCouyAmWUjR59y9Q3IwOCfGEhA0Vhz/d0Q0PouJl7pGdW0HboZO
MwxemVTKxamOOzP1/PgCZ42BOshd3SuJqODJyWgigTt95NmwEy0HmQgbDZwRov8f
f6X8/U1Ex8m3nIIk7bOkk/gpBH4fnfTsBhXoMJKw/PqO/qvSaYIOU+MrbgX4JJ9z
eyNjO3Alui3B1eHQJEFGd2+66M7l6GdWYMu6kvWFs8wL03nU8SyJUxpcGBYMLAvf
mqMiMOuRpGu9+Iyocucw0tP0cjMHZ1qLNBT3Xwz4Z1iStR463hkMSk9o1kwJuYu1
2bGM1xzJihT+MfcZ/ckft2YuszwiEGt5KZkypFArukkRzZ0DQ73atEE5s7OzJGvd
AHvBFpgowDGgDrC3zGYr3gDS8H2TfuU9SquYuqhiqkN92UaQ+1nnB8vLPIcmcxdl
uYtQ7eQ5NUupS1wZo7TEO53jbYw+WSoSQ+7drFz4VGr6+aQrHJmGngjRssPmevOn
wD2ad35Ow8oix82jaVJ20pAAyKPSocsIy+LMUeMh2ILEA5ZBKUfpuPWBgoHhh/s2
HGhAWzdO89aKKVpXcKTqWRqPk0pFQBWDe5qzXNo4mm6quGasabgiehOczQFrF44q
UWVGGKE8MyfPXKB1s83HNWPEusE6y5B6t8skx65BG/xV7nOd8/y99SXJopA4unHI
vrAodI7t0Cq4PRhwYIwCIvFzJQSaDIYTej/Hg65xBEcuBhY2hMVt+CJFgMMvHf/9
G7t2PcgCo53FukP2LqMvC0CKJwVLIwmrXuJn+YpZZT9WiPciqPp+Yn5RN7F9qFMt
MTAxHZDkLqTWbx+6vnMNpUAMZk1H6S1wvooVD20v/GjCqCXJh6T92H36dj4sSJDJ
5H61nbd3RBKduDD0tui2Rkbq5mOILCDMGugI0jv/8Grclhq5Feo6UWGlE5DoALmt
Uj59JaI7olnDqbYS405gOlPTk8rTaPNDfFWjulJUZNDhiztKx8XW9w/THh9k/7ze
eBncntC2Kte+ycIzwhw3XiMAblh6Cco1rgwt59pcaZw5Qe4VjYGhxA/NGeoBxBED
kFYEsfN57wXAQo4ouiWVPpgVc4VN2UlCVT2gYTdd57s3KTtOQpl3/inA8/+U6E0w
0PTSFsKxmdv+56Ko6h3Y58aL0Zpp3uHlBi05YThkhvRw8cSBfxSVnirlrBzWKNjH
9KMqxdfjG4KgQ6nGvmIh7NmMv8KKmcWHhBm6fYAcKM0yRMvnugn81e+lT8eD2d5K
P/9whBX5FYmac4srKdKdAWbmtVE5RDmZVpxXaPoIwMQiGuoN1M9omM164THIuLLB
BNWoCsD7bRzkh6TsZOoQDbGiW2U9mEgrf0HcSCr+TYLaC9HuDZjGL6QLbxd7ecSZ
k50l6jlTZVSosSv7PiUBK6aInmr4A+eKJk1/BdiZOg5pUYr8fRlCE3jXud2XpvJK
OswuPBJXRJ/7ZlSRZUlD4ZF4MGv0M1/nm0q9d5Km8sgixgh+IkBCrsOXM55SQf4A
7cX7bZEc30nt1G6u0LXFAzRQbDHbmcaVCjjYFQf3+B3qkGP2hounlSLygfyl8sBP
BgydLcLRnGm0SzklxBq7T9CyfRmb9Anujw5Nf3VGItqoC0Yfhcg1hcNLoDZcBoiM
8zZbQMQ8TDDaWo5vX2OaXJXCJlCSWYLq1bLuO89rQve2Vyq8KrFraiLzlH0i9Z0v
YWqf7Sp71GVAvSP1Dr7rUV82KU5vPI2UcbL0G1i8u39dmhGnun6GfESznsR44f0l
cix+jqfgN/R/TaKp2aDAj3EkFFsN+KKjyGAb7wWX7SbKimPZNNy7P+BzJ0X9uT1N
J4lXKXp4ODVv6nsz2QqZPrzfgLowkCSwLoVVkfBzSJ1cqQdDRYFUH/aQmYM+dPZ1
IGxTELq4yQlB/jE85zuQg+Llr6qrp3NtfpF9dUBiu03Iha3Oq752U77Lhvvbojjt
rO2YhkErR/c+Xxg+0IhuRmmSnLO2wmu0cee6On5VcTPoGs7lheQhHtt3+gRjzxhS
j27oJQiwixGjUyyXgxkmP5P641f+CgfOm4QeUpdQpn0huvM1GB4SeIYkmLjs6MNZ
sK4Fwp7a2i0sN6vCOXmAPqKVYOZLC/rd9/jt6oJJglrO+pKzJx74M1YRaKIHYN+p
POQq0GnhrmIJRLFq1fo27EN9YDB3SqqscacPyb4ghxin5yW8dMYRYtIxkUwc700l
ZGYuuzFmbeY1TXLR8OEWGz+sPDBb/TZETsD8UMvtShkVS8c+loeFUsZmNzUYisOq
D2+L+fn4duspi+K5CCtm+m7dN0tIHFS8ewaK4jUIKg4wETbGav8pelgac9/D2ncV
Sj9GgAyfbuNOpO870fJcJ+rRtBohh5a2pJY0ctlD2i+RyM6Kz6hWeHNsIOj5QboS
nQf7LEn+iXTk7DOd4NWnvVjzPHWeztKoo/eDnonLNpUnssn+HJoP++oJdaGmnXBk
srXfC2kwKkIsNA93o/8W7gYD2DlypZ/TqHzBZubtXQEa1Uh0Q7hcpmiNK3T97M2D
7bg8Gv0AsN3sQHBETqWa4KsqSD64uDcuNHWqnanB2B8bLFTW7RPGUrr+Xsg9bQSW
HrZw8vXxK7pP9klXPyK7J68DC+7AUeZ1lfLutQaKOhSSzX8sICvux8MsGX7HcPUC
hmjz32H4V4s35KXz2X9I4Ahcb9KP0HJ4dqeb5qkaZTbInVwjg9l24QVBOU2Vsapt
gFCH6SRHx45gd8nZbVZFzGeBoFJKr2pVQ2K0fYY+rSypwou1oLwbwqTB+BGw7Gkv
Y81j4KVDPTWp+OR8uZ4MNNC8lEo1sfIge3zsHNEJ6oEisRrBNWHZMZpf1jKWifhY
u71NebL9BZMg2p/ds2lXY7QT7dumb8rLZwl1UOwxa6p9dpuKsXSSPOYVtM4CulU1
AtG6QjIINeFwEFI/QmlCf4dbywDoBLQQtZI1Kr9j2UUZExh2uv+CZEwZXNGeX2Y4
R27xJH+UUivJedkTNZHtGOlJLFFIwT0So9OyltmDhNxZxWEcqEtsRxbGSz7XXfsf
yazFUoMdAeUq2jDBWGMQB0WMX3x5dbAlIJr+Juems9z3noMMmEbx8HAdYlpP4dGo
rrfuBcyMoVdCOL4cVrk9xJ3gT2T+93ukSi+Cwvy24HQevf+K3t8ZAEESze9luAGI
Ac4xGOq9+QO0FaA0msaNv7bNA74XN5Z6hFkDejIuAXvbktYHbZNUbLGQg2RLLIPY
zWCUNm8orQVFArsoaZZo1HJ6HqIGwNdcJKie/mVnFsun6cydLf7rar26f0l/Hx6i
lz7XA2dcgHOKEULKxmdv/+3A0HaW1NnqGjfOhqo8g0ksqxWR/JUo8akP99qGFuxT
q9hGGr1IJTjjzYc44CQUMuBoXMPBKjDl5HBijzLdzoTBJNunP1TFWuJeFoQvp92J
eVYWesWn51VN4eT9UggYOthWW568AtnCX4paozqZlg7icmepNfhW5ZHBExWp+L0/
fwHCP4QkY8xEJAqNHY1husKhbtw1HJ9wrQapOPoFTy9Adkmxrnz7VTMMSVUjKBp5
9ylEruW+oJDnPyi4lhjbrC/UAAHMgtpRRk3ebLahX+6VURhfZ6vAAGGBdUf/X6iZ
qLiZT8k2yBwcw4XvCtGZuwMYPTHwdBqdN14t/Nus39s5RwvlffrXlbEzz5S1J5tJ
v0udVD9V5KCzVvxYIL0M7yo9jETTEWRnTU91FxcEWI+3AgqFwhagliCtzQGEwRR2
rrGA4HNgZ7q3XMnBQ8J1J4eCQR+Bd3WLZQNOnEQRA45ekbe2Vu1mE/OV45oRbLc1
AO52pCeN8Pz8/CNjVJUmWxeg8E5VxE2jEwVDAiIimw+2/XYOzG1ERLf7zTyh06G9
6vD3VfvWVtRI/7UKVUHX+tbDRiMgjhPnm0R8VNm/1Y7vat2y6wU+XrfI1II5KKIb
IMpyLqq1y+9G6CcdPUXBpnvPV6wKE08DimDTULTR1YZEqJXvfxb3ovT4vXa+Tk6T
Vv7LntwgbLEHklfB6IWjQfT19EUCh3cNxeDrrqFml6/aAnlJnmA6Danl1vgJ62Gg
ntcvwcixXvKPNoa0BXh47ARBrvc6pZATNn0/YwZlVEanZCId9wl7g361StJtZ2lY
hQiyvC67b2MzpruB17cImDrq+LHy0Ma9Zdc1LOm6BgPcXEWLe6IsM7H9VCFOaEem
VX8ObEbKrPx3MQgArdi/dnQLs2aztZdyXP1IRWGYSDguSne8liI/Vw4NTJXn90+R
7Dti5S/p0vkAHDS5a32tJ/j4xzTBoEMgdMaS1kopafSOnv9h8NzwXYg/q0LaHzNl
TpmmA23MWB4L8BCh/468OVuJq1yj3lBi6QA6vm6OMYINMtXz0zwD89xhEo3YbGE0
1+jURe8vqIXsixSTNLZaxrNlZ6tvDwKepe0342wmeIMGKJji4j0LYYzowvTrmzBO
f3OvIo6oT2FMtA4kh/JT60zzuBvccY9IKd2rvuoD+QCzZbNGI+eSMikfBaMOr/S4
OM6Gt4EEW60L63tGq244ct4SQiQ2T7R5Ew9eIKV8MI+G/hR+zYTICIx4uYeSCWiT
McNbKF2whUaif9qCb0VDDaEFJMETFH1oc9J9Otr1K8o6pSY3vlnCK41+IkNTinsi
XtkggTGPms1mcbCaI1Xqq8CY3O8/OAnj7RHt+ELcN6uoOvwB5kG9ojF8r7UGCHU1
FCuuNPj5yLcfz6MsMaGJMOg0L7mudw/mgiVYpY6YGnBuunG+jpZ299WTryOoL7fI
wtp8Bt/AUFAoPO6H3Ae/NT1iGx9k3JkKXp9rZvE3MG5Y47cMinIQDRHgbVeDbiZ6
h2bLFH78EVOa9Dd960FREKipyMGVJaZSWaXHbtA1uZ9Yh1ML/JwHbZcJCshJoMB5
ynpgE3Id5M1fY5fI5DKosvc2xPHmW/ufwIfH2YiPVHNuToWISSCrtUD6XD9qNi3j
hmBVKo7nIuGq10sS3g2WCchjYDlUwWzRmAQLNw2D+HeBiFphb4QdZmPNTmhOrOCH
FpObqG5jX71e6PUfCcs7a6fJYHleQVJ+aUOQPfe/bA3NUquDTJzIM+lzHnF1OZsj
3yzz20Uwoo1BV6s+PFtxoDBTC4g2tEhi3g6m8lm3wFamw+H9LnKr4Ui7pwLpSvkB
xHoql422BoKQtPin/nHedF60ed4Z360Ejz3ZSdy05kYYowZWPJz/xF8krupI9hbW
ShfuPXysDKH91H+FFdchgKQkuiJoeCvK9UWc24VlCg3D+0slRpOa7GkavN7aG2+A
vUr4EEo651pQCkXuAXRlKJ+QpCa9lWGSWa6MmZgtzq/JatvZYlzwzWfiez7/YpRd
KioeCpyFMFAiPzKCLv8GdQRuj1iFfFcMggeoK2yiOkBtWQHS8remyOhcqzoHjrYQ
fN89QodogmieVRF1YqOa5p59fvGyh78aUZli0z5JWilf97W04s1WRv7Q7DpTkf8N
TaFr8LZfZh8bzwCEh6cc0G7DL04anll1uLfdKubpvjkTCQzrCxgmPaErFdhDDnM8
BpRz39IMx/6QN2dLsuiZGF2k1KSaf0oshqXkRwZqLM+cktALVoak2XgK0Luj2VoH
xCRcCFnUBqUfGbQXra03qY7wqKCpSaJy7vwX6WUCRFbIlc6e/Z1bSx37polPSQ4M
ovsmqG7vcGnpfkHoYdG/6iOTwmtnQxps3z574C7vRX7WJZLYx96rdoBR+QdCTmIB
v8x3iZkWhtZ1rz0fUVWPAvOOplzq55IMmTIEzYlXGtxJ6BQZvjFVROba+3zM+PIL
FjmSfpdYYbsJbOfScozWge1VXWM5kjF8y3VpmGK2Zws/ojawxWF9sfqtQiM4vZFz
HmeB9+Lp90GEO9oWi0R9vOmt1EZgys1ByLmujCW3vYhjIFfiYc5sqztTvElMyf1C
DiFj07Y9jCIRDCj9Iv+T+t4bruoXQPbTzavWR8dH9ZkMdj/ygupmwspC8wMwWwrr
VWKbk6eHYgLSR/LdsOsLkfUmGhT1MjFNvOfgE/9BauniJ4PlJH2Wy/Chjtbo3zy4
u0ghSZECpT1QQzQtWsi9POhESX+BTcBZfPUj/2Etb40O3ToswcPMr210AN9uDmxB
iihoTCfs1M95s/0q8VSmgHQZLgZWxHkp+NtyDOx72A1H1KWff70XuAJborOlTH/l
oZVTqcHH0jQ/pRSx9pBHEol/FPlgTQswRoD6bu+bS21ufZc9XLEse/WjEU8yBnPk
pdzx6MDXGqWQjv4t5PdKMV7LAB5feCt19+W1+XVoNGXK7DqYdg+ne84eehyndFml
ync8N8CEeduoQdOHj4QFsyhxjWRuFP8E7hB+kM14SzlnFUL8W3OhtMcii8ELA3Dd
Dgdp46GU4zXrdRTDL1MdZju/R7H0OIkr1ZHq17fgMwZciIrTEZotaVYqzsvlqTfp
gnTm7uuoyxPJbusN8pxEFGMBByMKZLKXwHcphhT0Tt1f5ZgOBGUED+OQQQ1Tm5cx
HChR8du2drk4PHtzrEJ0CiIyxsjjf1un67KbdFD58lOTWZ/jh81UcIdlGCjFZ2gl
VU2lFKhKGirftLFpAjcPEPg2Oc38VcXjBzePfN2VcjJxcYeiCeCdzfBK1ib733Or
HqIyNiooU8jVns+hkZTmWSRwvPqqxTDl6+IUZEZjPr2T3Li4/jle4sTHEFC7oTSN
hpnkPlqZ/6FKAsJ3/SfUWZSId1PDyMXonPOeJZvvXhRL1oTq37Oa2gJZkC6vl71C
VXjD9/wYBdEW8YIeu8m9Hdas2USNkBlqqrida9FS0TOW0tauexLtJSZHz0yzHZ4R
jTJDGppMUre5Kb/nqZdI4mzA0dNDXG9I/ubbxQiUNvt6+EQTyDw60BVD647llix/
Vf6wc8QQd+P3DBfKF6wrri9nGA5mUm4nA0fsmySSQm4tS4uhQN6QAXtMqEpt70bL
LrVL0INVE/in+j3t+AfmH+DU3Uvjapo4OqUnRcaEKty7OT/EGppB23uXg8/1j3m8
v/IpheJcm9FaxEACQIOnFQtrInpumn7TSSQ43rFB7kmi4vpvo6P1e1qBSvR8qCji
VPdFUMdcd9lPwbFj6/TgnxQGWBb9fQQJ1p3zcy+HWBNr8OEDndo6s2Oz3x5cf6dV
wwj51aKaOHB9VgQ0n8F9t6ayu03aP7Z6F+Hny8apiIe3jY0AtC0Ji4fbFxpaNi30
qWNlszQ1/koLitKYGe1HDDPeSE+FDNYql0Jb+tzuv6dPavqqv6uqwmVDL8159hl6
3Lpc2dvSoZQyJKGzgcZhrw+dZqkZZuwPV7US1nsKwMmnkcF45pKnqDtCnzGXt6Rf
/f8hiE8lArEWY6Zo2td4kEPJdMUS1Rz/9F9Kl19TK0BlKlHGwrSigRotwxelEapP
UVerXzOmztCSjlC1hGEHlrwJG/2MVGS8o7sWCtaZgHU/i71tfXOcZackdaS/qKv4
Zs9ZiBIR+icLpmNo5tEEQj+1XmfF0AB8HyBoc7AzHCc0PtSeYlVN5rFdFoqzmvMD
IxaNGexqr/bKxXkNpyRcrga9iPvzveT6/5hV4SiOkkc=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
XKI5m1KKLQ+3RCK10Lsge2uoY3LfaOI0hDeOtlchLhXW8P68V9fwqs3ELDzxvv5D
IlC7GTgYqB6Z+vO0sBQQ5eUSiY6EnpSzkLhPVECFXuP3jbDrkteHxTaWXKimY4TS
pSC92RxRE6TztyXFFEi+Ak0GN9X2Z1v+7H1KxsXKDXs8mseg+QK3THyyluyySByw
j/8HAAXF6L3ipXHmlvufexvJ1PJw8GWkHVh7YHmWHn2isMwzuwptOI/gVkbXE7Vk
rCagLvPUv0vG2o7wfJ0pFzCsEl0rLEm+Cv10pzEY0XzYB6TPTM2cNgJe1DlCzj6o
mc2lBbP9RyxeyVvFNHcFwA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2000 )
`pragma protect data_block
hqL+01lfRww4jil1zuJEGKA2CJFH+L2K0xLg/4if7Boo148oWV1JuCkMdTX6umVl
FYa3hG7f05idWanxAY/QlmWSDgaWQGpInMchamvn3LGZqtcrWopWLliMQ69wV5P5
vsAJGGmygnwnxzgN9XuVdwS14yYfGEsIZTybICthucjexNj8URS6A4e6CLIAJAM8
LiIpp6/Z/wiPPT/vM/161xNTaK2cDOLVl/LKD+GweChQDIW2qoyacxKoF27+Djfh
cjN1VPt3+ypfYEswXY7jkyUH/SgRwawfXiqRkrSXIyL4XuQEmGyG1GQRKqQ+GBVL
quLKFae3o/YFiLKVxQLYPpR7LDVwHPtBEpoZL9jB//At7KXP7W67NDZ4ilbiStq9
wU1H+okHo8Qz6rKriDB2L4IUZvFGgd2dTWyTMefCT80LVrOCUpaD+wDuvtmS1IKF
dWPBVZQAMxqKQ3aMIOCFzA0OGzByFNYYVGdUDhGrSonyB0CF5jp3rhbOGiS1syJ3
nsMYbGazCHKDgz5oYpo2brAqXFO8PQN9WDzvfMsR6D+FioBlg3LSANVHeEuLumZ7
Ykg5yyQf1W6tbyyQvuvftJBzB/ds2zUXBhK8ijtrQ3As1h4WMljkeBohInfYP9Cw
NWGmvzqaYjZlWLuEZohL4dyefFIkfc3zQV1EtqVtvU/k5ijQ63R+0JSJhqhl45fD
siTaLspXHxAKckjWdxADXH7tHfoxXMxl5t09dzZ+Pt4XCyjIV4uyg1tHj5bw9SiB
b18kg5UnvYZw3gdFuDjb8DMxEC8PcPZhuvVU98Zr+GsMlmbR2zZxPUb/c60nosjz
Dc/1OlFhLtXdv7ryEQZDALuxaQV1EBb37eBc4pD066Xd7rlf4d3RtwEAhq2TR7K+
NfQqiWWhHlrb++z3PiA+gHYsN3TgSolmcaXgiOt373QXa5pHn9iYn2xRsVZpP6ux
zOhIf7BIdCGau6RJ+b8YFrtvQg/gEV6OeQ45BFPKVahfGMtmeV/geNsUi+OE/Qbs
KePwvQQm0vszfL/ZRkPeG07cUVpMjGr0s52Iqm/mSG1MUkzB6V4hnpf6kveNzviL
6PypgRSBHzGlo5wJyQKpo61yKuKzWb4GY3w8o33CKnpVFflJEuLyZPasaHWs37do
5YKkJZkQh/jBxSScJ4T5rIaQENt4pYyZuGQXTGoRgk7emRCqb/qHpRkD46NQzELe
45gQUPjFCsapHgXlkzLVMQAHC/k/iz485dE5S22qW28TyHE68wA7AhIfEmUhMrSN
0l6bl1sN5f/MRdau+2k7eweu3GFzjSPpXdWpkJdrJrOPlx90mlYj/PK1mz8zNUFj
KmykvxdWnwxDAcsNLNnZ3Ipr7ON2aytncdadm1xSUHbww/2wc4ZNQNMjZdd41cmp
Ikqps9PZEd6BrgY+6WLXGmNQuYp/M0nuLLbuujx0Rf2LKH2hl3nRY+6XEaEFXIgc
BLvr8iEN2j2iFWK6XOl2fxlSvDDiL257m3hzy1iGT7R22Ur9XikkTes/lhVrdllc
FVtdC0JSYi2HyDhGkA8vglgfNTKmeJI6NmKWiuHmUguHesdztX1OqEx3mEeZOHAt
3P0cSJGj9biDq1yY0rKraVEbz6C4TYN+XZZS+4XYdUxdpgJ3y2a7UYW5utuUF7DO
z4rHGV6X52O4tw1I6hYzyQAQ7yMUWaweZ9JQTn2VxywkcCuID0g2/LjbFJbRZMwS
kyYlSS2VYfCtCTKWpu92c5zxkuDnsAqTIxIWlqJmrmqlpTpxL6ZH5OGy7HF0DdRv
8olbMVT0Ino8YNYQhBCWVg+EaNtS11iaTsS9n6iHPApK2dVJ5DKAPKZCvJ8DfR0z
FAr8HkWYkt9ylXfHa4H1u8jQWNZlXsyCkeqUpgUCf3YuZ7hCkN1MNSy1gKVH7Izn
qa2z56kOIR63RDV3BXgCSVkweCVK1wOnAI8Rm0JRWm1gjbFziHEcYmxFKB7Hb+Ad
vyNM7lq3B8EC6bkbeA03DAklUpSXBNdu7/2+pnbbkOT3ClV6UZpySIcx92bl75MA
z221M2edPctqzxrmcVQx8uNEmtLSVnhwI8ZshPYFHEfu/FTaBuI6CUHRx33J37dA
eYe+qZqX/cEax9qG/BVEORG2CwxNfhTDi9q2pTNozMbfZqWa22EkBBIiB9tqC+YZ
SkQtgKTusQd2yefRUf6PgX27CW/ETJP1U2gMdrtn+sgCqzNwdWwe6zcj/oh4uwnc
sPqfxF96yo7kR2FVGCFvu6CI/fTTWEMgtIR8uFjfpe059huBPIsalsx1NeCc0/Ze
Tf96ekEFd118hHClpWdwahYweWT+q0Vdb+tkbQksuJ/7Wx+oqFmlXAnKGCRsLxM1
Of9mxStmpVLwCk8ygBR748TNVt9smQTEcRWxYm99NPNctTauHUjyiVuRghE9J+/V
LruAKGoT4OotDWDVjk/S0IIWakpbonhgJeiK9jhM0/20g87WRTAANLEWEWKRChV6
sHoIpsRc63AZ86+DQMmeaFpwtpUsEpynAlITAbVbB8QSUY3Jei7dOo1u/CDIBubg
+W+gCizYXpDeLfzxcCpdeL+g/JaWX6DNm2mKudD5gCP9EDriqrjjjkEV2MKgpEOK
0hLRj/J4RgRuSVbXxw/LvpusYEXnBPvr9Nf4ZEbT5jo=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VJixlraPrIxZBO8nO5zQBFXvzNNzivd5EBQnniKOinjIZnAYieMXbQA5F1R9ABbT
44pBXV+MrBXHIEpRlpTXBOeZuMQKpG3RRE0hzuNOHT8q+383/VkEawtcXU/MxAm1
B/JBU1gw2YOygddPhdUwF0VEKkHHiuUubVPW2ZRHtllmUXvgQpUoQBPohVl5Y8Z3
jnnKKrGHLzID4lfv614tmJTIn+iP2LZhxIbDN6/QuQyNwkEe7iecDr7ESEWJpkTe
3s9EfCa6lFR+rRaHgBDxWn1GH/4vKzBcxf0AbEGbjtjuF+UlfkwrG0azT8D0iK9Z
rQdoyO2WgMRCXsWuiffv8A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 22480 )
`pragma protect data_block
M8BqAwK3nSgdl6O5FyyYszGXsC/07fH5wC5UHejS0FqJisjqm0DExRDwebQOwDdN
a8QVPGzKwj09sikeysuZOZ0Owlu851wQ3gPCdoH4FEMpxlLbj7YGDd5nGxgJGvAE
Dbep8e7Qr0G2Zo4EbDbaJf5RQ7fowjuMNy7zda32CshXbGb25qJVUVABC1vByOEf
EDd1NsIfItrCBu21nc8uaecG19jhxk6TnohRn9eJlEQIyr1iFMrnLv1zUoBo+HCV
8+hBlqKGwwaHGB9DTnaHjg1OEX8EhhmfGx2EkKSPOHEykHbAsJjuB5QCZWKYLVAB
k8iZVSwfh09qTEj30N16q/fQfEtj+FpCSKUZy6Gv1mVGxQyCeVio3ZgsL6yqoTaQ
XDyjoodUucND/U7e4KXxRbVVZDGy0S++Q3LLPjnFEgdoNGlFCSytmxN2Di0N5fKv
bTZwsfKLx0wK93zencS3qi+RlHrQ8TYSrVBemKSoiSTFKQ31mVLR0CRi7nF+W6NU
eoyzj3WtzGsIAW04/luQJh79HFYuKPngkZfQZWtSqHBRfStry1c33cpLhYQs8UIv
XIxy7KtZHDyZu5nF1JyXTSTJ9EBRzZ4NotCc1vKeiJYzTFUCTCuZrUiDOCV2m+fX
l3YB3sawc7MOl/zYclpQBQFPvmJ5wYp8SdEysBvRAw+FoB3NNDbVTIAFeQrZv1yG
zbYvbtEiuux0nS/28z+JlH+yoG0K8cdPO7YCU6YvkUXq0BfHrwjE/ck+R1Oh/R9x
S9XTuaJu/0XtJIwZQV3/c1ZikgCDmjUhAvR/80NUuxhsMgS9ojlD5K7Y2T/Nm9BM
hpR7Y7cohk72h5irJzsM+sBuQHw9J4GHqvVguVEsODmFu+d8JD94kHHUgcOgA6Vt
uG85n9udxRts4Kt3TP0tExyflW8dwQO1fTzOiUpqrl2f8e1h8yhvgawwVBXzwk60
wNqFxwoynGMP4iYoA0JSEkrirZfG/kp1OweEmH8Xkk9aQ7Eklhu/BdPYVS2eQh8P
FLuoi+6BPER55RaY05K5WyTb9BqMGT/Om54nIz0HjfvPgz97zBd59ugCWkPxcf5o
QN5twMNsxPhYCQYuqrCnGse7QAZMRTSTEalfu0CEwek4GSEOMp0+eIz0bYXWOUZu
a42yte1oBpFFPF7JVckPj2BysT6THVy9SGo4iUfiOkGCOzHKrrj9ygRz3kXr3ntj
tvptrWGVb4z+JG4cUbnO23G/0BbgpEe6dvCuAgUwbBfKLQHbQvHErwRKmhPmYm/u
JbSLGmKx6a/2ULgpyzLiiadi9ZiL8h7CrUn8MpXH+1QHOfXYvTEJntqIrhfL//eM
xvw3qDbhkMZyJ4TmuNFn3N1jUawaUJay/akCAobXnkZ2jutCJHkvo6jo1NNMXip5
xuV1IXrhbFjwRO3wREM1DX4aSDI9WtvMKZNmORfzOtlYXthmqvPvKnLHjm1LRmqj
3EPNsb2+UM5faJRUpYt0g21FbQ1UoocP4jOL52QBY0T6zwOfUNNSeqch+/WmRt8D
ARXtONW12JyT8rkkDDmdh796Br2eHr6m1zOSbJ6iIswre8KzsY7R9ZMTLmb/PUPa
fDbp6s1XrbZUyCBCQYU/r4BpCqQkwPZYWt8Pr+l26SEIcnWJIVv9XbFARoPaeAWq
Cj2OYgA/m7eFw6MRgMYGvJNbKjExrJMl+7TPmaMeoimkscZikxR0CjJKv3J9KYhG
fBl/WlNsn3Yf8Kz4APii4waR8GJQ/DukFp6ajRuwwf7U+U9lW6lCUuVBqusz7JjB
j0f6uNESKpVcl7W/Z0itC3np+Dyqs1zXAItf3Wl5k1slqHfbchyAkyd24folv8GK
lRIMrSb8QMhFkpudEBzBtTEtqDMKtHKMp4se0SClOU6LEhtRqVImGrzarwlogoNC
9WCiC2iWYCYIWpwzebaxICgKqjHNvRXU2J25Yi6n/wBQ6mdjFT6lhrI3CWD4zAfc
pIyHwpXlqZFbuIPsdc2+a+Ca/uFgF64qNcktbxaPSWlDVwjHESYdPIKvn5s28Z5c
7oZ8MXE3hE1AAU+XGWoGGh3vKJvtkzs17RI1Ge06NY9jXLP2B9egGZYKIpF18AMH
cGktMad/i6mQoV/pTSbC5VZu+zlHWZdhjKbk4n9udaEgZSGrnVyWirCJ7b0GjWdZ
TYDKrg79mdWoiejZ1UhIEI2lPrfsrfY2iJGM8BPlqTk8XO1+zkku4LE79EU4tNpt
hL9daq/f3u8aEILoiSoygjRjjKlZivKU+2v/ShCsKXlzT2QcqH68h428qeomZtbA
RSF/eY81BnNrkp/RjdEB9GEKsYA1UsFBhJZrvNvpQqroraqh7engHJyD24F6r/+d
aIZ0Vo/ZRbuFbwPAmCCbY+2g8gxjNnr5eeuLT/890krvEqU6qDosU+a7nNF4axVf
5+V1IyNy0T0w1zLksomcVi4EDlfwDjq7QratrKvmSQAT0RSd2g8TxxuBzOtBc86v
CalvLfBFiWd2FZI2DYyFbl/PkUtR15pd15uzRv9j84gx6P0553Zkbr4GGBfAWgOo
AXMBFnDvgIvcQcO68Ybw26VjxaCmM1MnUm3etZjEr/AcyJPD4M/SagEfVSVswbVz
x20vwCHjgr90LeumCdpEKTpg6eifpGKgfI3q8wydQVSIeT2twA7LxYEwZEuTrrwy
/5ck3+F9KyuQQYgCSuFjmqF8KSlSFFWjv8MIiE8mKfxP+sxAOv9qJmOQWtoq5Bkc
IzBJMq4R6Zv8YPfVtU9bbeEPuqAWoQE0a93qyNtSw3GZ2godj6lF9m/4bdzhsfRQ
rxIi/euChsD4FMKeQ3J6hhhhtuMaV7f31ITPsKpUHedsi9k5ZxH8ft0B8WVkj7Xs
IXc1x8Lp3y6IVqaHMgprXEvN2oGAeaiPpW5GKtpQRC8O1V3W5+ifUAaX+tkmvnvA
0fsUxue1ey9GsEBvnwyvrCxwLFcTWIaLRYo8PP1Km6Vs1ZgdaqpZigy2row/CmXg
3CUIsUHZ+svmiuvHChBtVUtXxpcJKty6Fyr1qjFdGu3bgL3HePZius4TAXhO2c5K
zZdpnOsHij/jK2jvPWpv6xCiy7r8XHU2Kj1j2zWvDlnE8CYYNg7QVPas1fH8wMZm
jiiFHk/EyTc9M7T7Yd7YuUIr5MVJr8syFJyvWctXvhrvqt3FeEr/VxAV6e8/GcW7
994Glk55ZhktsMBAKAzrMBMoJGYAupXH13xu6Ege4br7Dj+WnbTD6Xku407GEaxt
H64UDH3fN1QKGZRbnyZtygVuW1SN5/mr0mPl1BpSY3LAUfmrlGIJO3Yas7EJsnqG
4YVEjLhpJE+hsdOlPWb450t5XR85sDgxCyXvzB37uijM83Q22vCTbpz2ky6MZlyD
M5qNGmS2o/Q1t6uBbo7Io4PmI+4Y9K/IjtynRJlm7UQKwyc2cqlCq981qPCxtAwo
AmSSnTccDn4xifc7aFktK/hA0kBELL7yk16VCwkAYGyGvT2n1mg1Zvtzo1Xtd44Q
dYdNuKDOaq9pU/ETjKTcTgpfx9aW/0Rm4e6fdityA3qXeACVrWPkCd2mZ6dfmU4c
JapKkMTgKl6ii9+AgZ7lRXsoQnnJutkyAX6eKVsU37hp5cWh6aE9truc8VEQnRi/
UNDRrlcut4ZcCBiuyW2GlXvx94srybxWnZ/842KOK9YhWgpS0JpjDp/9liou/J9q
64Oq42/rF6gcJlnhHJgVsDAm2jja9qxhcl1PmEZhC47rrhLBhGwcCDvgLXrAvBoQ
0dATkUog1eLF+58GGzck4uy2CwzrgRNffnfwGmdvxfmkCM6kwbvvDpHKqn2lILG4
KwTs8nL/oW+QouyuI/8FwQbvbHnG0C3G0PXCeMDKf9DDkTNq4YQ0MlN7Ay16ZXHA
AjWc0g8LRk1A+GmXHMY6/s08uLfZLFZx/Bf9q0pWG0J1wlukpmhcY6McB0REgsBV
jhVWfdJUN35SKsDCHpTpBQ6TQh6hFgVHL7l+MApxqzxIsxfGoEs20amX/1xzrgTY
miNP94iJ//i/5frWvdxqynAQZ7mpx0eu5o6AUc+mwyAtx+516qDCKtwDEJzJxLw2
U3m+lUbldjqBvMsnBit4mF42RFIyYZOpWXt3W3ZfvFf2deBulg/nAL9F2kgVb1Gc
6R5ENu0YpEroPmiqgRBenzAndw8FeTRNSY+EbDEOhpCush12RPTaRFEhet/RmlEl
HXvJliSccTQPd4eF2Rkw7gW+dpsGoYzr/zwJdOTk/LWplZ6W70xaTkQwC3n796ks
SDyRp0/oc/AX24vZAX4uDUnty3NvS6QTzSnICPt9J4rylbFjxrXlz/z3T4lASqqd
7mv6GvjvSHimLJHLrkp6VbCxasHktbNYTBu12i2v051anlsY+GxZwihZqxDe6GUE
fNvpdEY0V/OEL+u/rbbEC6SBnwzAGgoXFP6iDLsTcLVDAVvnzWveuKnnSVzIvmVd
ridv9ZxIaAGkRnEg3g+3a3mNsmWMi4tM8A8LkzbV+h6YAYuyzWyuFNtO/038Yx80
h6XOhi5znJ7KeXqmhX+uPz+TSPSXiFfyHnji5e5Ihb0CVv05eG74Lm/M4YTg2yIk
IBf1l7qCJINKSW+TbdU9FEgEe5Z/AvUl7oBM8AOhuquHTCNZ2chzhkNEBhpq0pKJ
cAHshxOxY3LJ7k26GAuGfYzOPS09uDIioctdBaWbevIFfZClmBN1P1myWASzKxxP
I53cEnW44U6naMAor3dmLAkHA1K/kfBds+pUlMMzk697QznN26OhxxpePQPX7Qha
0YxotD/yX0rxlmiJjZILO3w9VTwqgddATqVpNZIppJfK4pOFusJTvXFLN/P6tN6k
YuFvnf69bksXhmzMPDv/yArus9p6rcMj7Rr86r56DRIbnTHDcZzesx1OSZU5JcFD
s9pv/rxYrU+P82ZNCn0OVh6KMWQKtyOOkbweBsC9zSxzhFBJsfxThOq5KtO9GaPv
euubU8E3EH9OYm1gf6TO3MuWqcmItSWkI5dmtYdtPZcyu9fR79hf07f4TGMtUhDy
hJmx3bMWDVDb9rUYYTeFUYadjsAndLaojYmQ6snPBdwC1V1H6/2pu4R7zpwesg+T
R8vi14xkOtZ5vxBfBnC9wqnE67iZnS28R0tOccwSzqnuZX9dyJTUkTn1rfWJ8IfX
riiiH7kKu8T/XpMSgramU6QskbR40cEqmeOybecxifzD+gZo9FK4TJR5X/QdBRSm
8X1DLv3QqO2SBr1WsLV1V1zD1qRsPPlBrRMT1Z+hiumBncWJNunjP+IXnaaMtnlh
KpABsBhC7pOMLFWzHzmsHcWwHm9S52y5JhbYE7bmBn4ZkJbAoHGJz/jcKpQhA1rj
nYwoOxEb+CC5PQ9Leo3Es4l8h3T69u1onZqegeTfWMyGGdggwUIwvv1K9qXZ64ZI
kxKnyjoCBbLhEHsBFEn40C4pSCnW0dRHXySrP251BsKsEOWHBPPjMKmfDbHMM0Fs
DiROHmK8g/of9+UMjcbz81ztneYbiAWWc7vHv/F87zHtMXgyf6sRVG/SEu888zC6
yCUTTa/rzF3xYDJ8JVcQIUj+fZ9k18eqOvcEK0Nn+FOb+bxmmD3eG+KvkNTZU8a2
Dg8lBWBoblnqgwV1ff94nAL63Z7Hsvti/NREOD3GmucSgj3fJpZh4JvopGsK0oh2
mEq3K2D8qFYaIQt2zU7HwS5gg0EnXwRWFoJFb/o+UuEoUH/8dU48Mhla3OVyRytz
1WgkGmPUm6apfn99OT3O1dMOG+Gqx1N0BOvxzdsBXxgCON39JTdlznY8UY4mXSxO
HCAHAaaGNaukRYHVURG2Isefxis2V/qjvyY2zabzslMriJ2fwhUiiPryHLYi8nnm
PoXg008mLdAOHMtLEQUeXwqf81uwe3vVDYKXtPsEd9GaXIPvPwcODTpc8kFcEhy+
F6TGCF1is0Jej57O62X6SeNlkSb2oAvrXyXwOtnID3OnNufg6HLyyz62UIefCwHC
jcqV7TKmUKV3WlcZI76/QUDwlu/AaIyiZF2MLBusYZoV095NSQuZq4/yhbHAO+Tq
h5ZoAC8oCfHILx3jEzh7sAMOWBhODHLR34GVm79Aft2802tPpE4/sNUqgp0oiWxv
o3zXxohfsEVJITDNnw/BN9OcOHaL4YWppCdfMH1P8KsI4heUcBiP9FtSwtjJ4NA3
47CLJaD5Ztk2IkIr0LZt4danjVDLqBZAQLasHWsCUY+8TdKeBXhL6rMUxG6EF/oD
5JM7iMsi4sPwBv5RQ9CWSBQcPwIzipLKeNcvJCJmNSNYKyuG6npRZohBOq+4Xx7m
dtilK9qh8O+uZZ1Bh0Q59NtGSXNp9OPgsLpzigoYdE2hXRyqdgVljX2YgshrDwZE
PcujDD/fP9/+ezg24rrx770L9ElXYtQjf1/LKQDmKYDvm+Sy8ux3YxCgggoMuRd+
+XXw/+LvKBC5/iz2RgH2IXB8NnxkMz0DxCH2GCRL8GMUXycnIhXbHDP7H64bw4yB
VqmcjJfrkcp2ECWFyKkugCyC0+Jc1mrSS5OgWj7wRtUQ1426i7wQQ5ORa6m61VwG
oIWu/v9H/DTsrBwm7q+dVoWk3nUhj+rHEeso0RmEG9d4S7wt/6VmpLQ60dqFD/Zm
zwxJ1FOc+n55ypuGRN9sZgQZUqbZvFu898EoRpzohnI/9QWP5CaQkDKF3M1cP3nw
7fnMiaLHMhlXm/4uZX+62zMEb05Yw7QeHYh5Sy+9iPQ0dokkkFrNeFmW7O2UtHh0
DkRpSt6fT6uirZ+AxApQ/ZmWGjXmZXHQ0hfeFmbG6h9RHQzQsKvwDpaAWv3ltoxf
w5QNiP+UT6dB4rb0fV0nZDQWkJEpRJ0ZTkL9XCeSFhPFEpd6oDXwlQfJyDq11LQc
cDlVLtvhSjvPt2lVqcs8tkqahMQgOFeXJW6eXgqw/ux+NvS5uVKgdNQ3eBWDEa/e
Xb54OIqOGHoBiWpr+887H8zW+ZkydoAzttDYeuNneur6CeVzVW5GIJIUEnFweW1v
r9+ZOY2iwgcumZKI7Y7MWDI3P/1f6fNM1t4cIWFFmjJ+g8TmcVvz3ybw4jH0Zkmn
yEMUWvQrcxotURFmxmvrhDVEQ2jJ5s678H+4B/R8xTx/iwg+JizRHu9Y9KlAUAdw
D1jhbF8eigG0AwKn7nXtapYcWEHwN5XncgsID8U96Pik2QybKkDYMzoZpUprXPR4
nFzRyiJorE73AEJifWYnrMQF00l+6++/A+3wWsGK8PAsXYhRXA3hwj0pSS91QW8o
UilEenF93KCrHoisYBhGHNm/GC3JcmlMinNhm6a5sQgFoWr7YM12DHsb3wW+P9YU
/zz6xFbxBpyTySr1U81DLoYQtBn3e9TkSGBqL+2C5p24KJPcv8MItQPfVY/JBwYV
WVY8nRPmhAKauN7hdsaO3UWRKesv7Aj2bLWJJDGbMN6QnV0aXH7XQkYlGQELgInk
glASnHRcqYUHxOTI9QpbppdKdCExMgTdZOKqGYMSN2pGM31u/Fxltf74aa9lRUsY
6UuhBVMAK0uhkEnTVkCL0Jx0tXUmIMIbqKoQcVOhXRgLDX+rtbXsihbsJ/M6mVlf
VPLUwEhCGNC3e5pCJQLMWHZjdnzm/HzjtLuF6GXtwSi7C3lKtfM+nwLK4Hi3jR2Q
/lCxvj2AezMgLiGq2pJqBLsjOs1Q8a76t1rdjD+mEOPOWVePZhdgZ3EESC9UTd9E
XuS6W/3XS+jmgeK3Q5CoNJ1hkwYewPoK3XVZeMdbGP/if9IpK66DMVVVUaHrSy/t
WvxxLfmTpGJ35Jb0uA7yaX9Rvzfcjb9nFk6ZJ38dr4AS1FD8VC/RIUKI6FbvSJ5b
ZzTKQ3sbIlWU/U//hClYeJhU74f4JJL8WjcvAI9J8pf4hhiN0lIjJVfavLK70wgX
l4l444x8Yho8WS7nXKQF1rW0ujh0DZFTmJO1cQ2TAv89JLjqy859UJYM7z8IEUk/
rpSUQ6LVJfbbHo+4MAADe3NWd4FWRdlNyV1zLO8M8pItkPSdllQ7NIOkxb+zwG8B
k9Xj9OFvhHxhHXsHaW6denQStAUqfWfB2Qbsx5SaCzAJWUq+RoYIkh+D5i/bQD0k
Q/pygfYMyfse98vBAtxpHteqqMFoigCjeyIL3JHaepGMSFP3emLrrUX/GshHO+Ex
MwP6MAwBv0rqRWYPH5Q62qIvgRtK3B4dI9MBz6IB9fJw9f+6+nnjj4fqsGeruQsQ
FS50opfOFJl/IkldkQxbgnhLBJr0fzskyIN2PzCLiy+/15J4qtkg7scRQvJtZ1Kk
HDuk+emhBgwj8ET/RMF9oVJwksaLTJ3P21B4/Ba4nqmSl8SISsOdmpDu9OZtMRbQ
wokHo9b69dME8BXyYabnZeZmjGyIq2yuXVRVwD/eSk9BqQK2LzH9+7WErdGAZaoY
E2JFICL6Ng6NHU49PzDP/Ar9sajnA4/qI2iZMTFH2kO1F9wmrfvQRm/0PmOfdM1a
uTmq2iYzOP2yyyjj5AN+bBcldrdbkOYHFXzTVN4GT+Kfg9/D5dieC3JsFQbWFbMO
qMpMuDhlrxikgjA5WWmpNsC4JuGAPEmoQiiWACHhnMdmLV5aevDbL2RwHmQBgzLq
5xDeqJsLFbyq3tfExwHVdSrD14q0eSG3DS6eGwhzqNKmJwcr/hweZSx+hBlJxbnF
nwM/Emau6lJOlcqXKcf5ATnGcEnLQFkfcNYQDFSQF+wOUdtOQ16HCV3XIJk/Hk0S
IgreoPlT+enba80nvwoj2vkc2uT1DkUQv87SPMDa8D+E+b+K7jVucz0YaO3r7NP9
kcGaRtV8bvqFTe69mUrVWB7AbOXfV13SxOf2UPl4+7Iu1GRouhGW508OGOZN/s2Q
zvSy6Bm3pXANGo3Jk4ndkakaR0diRoT94rLX4rzmIAqkO4A+inBXTEGy3/L573DH
XShO8QPtaOtsNLRKP1ChHUPdGdZ3dur/2fBhS7n/6Yadf9eI8Kw2LqEtLDUqFkUV
s0Fw7nF9ECAQDubbU+TwDMA7Ep9RpGccGiFI8/0ki7ws/Tnxpr0ZOwNzLMuq3oPf
xKgKoZ7XHJuX5thGGxZkXskjdhZfYfoVZsvMPH870MmYQDMHFH3kpXHeCuY18Y0z
6FeyC6BfhCHyiO47CxTuquE8M7A7rtl6fA0n/slIb7VfBOc1vE84RkFKWkfiBGDc
+tagzXmpajKWOihFsi1yCN0Mq1qtGF5FmEWNc768JcC1QHP5hG2qXIWgDSLcaI0n
yBGe8fW6Z9a5YdBCeXYr+1LcJMW1/GfPV4zPVqpW063wIpYkXmofNgMfY3K4MNFD
ZnUirG1odObxqL1ienjYKDbUhjt65nIfNe0q2AuVOdzfdKL/sa/IhnujCWa1L4PJ
EMCfBH8h49GNyAg9ptgHhuUpBcaTtg7pKkibO+vWsXjqmbftiCelxQZhYzKlJvB+
1YQkQ4SSjt7JPqeonYndfEeZAchhOhEpNDRQmjo0CJHtY9U5IJkMS6a1b4lEi2dC
Z5q8eYSZMd4RBtev/17RWV+zGaqAqVxHR6CLWE8p8jdfYk9Xi6uHM9YRsq/Wk/iD
tzuCf5NYUMqvM6L+hQwmxy8p4n9ohQaDek2kOO2BPwzZGUSQgJLs8REEh2ZP8jQP
xRN94m7VlxLLzsTDzV1p6uTR8Rd2TtPDheVXnKzaa3fvGSSV07/uPf9+rEg/DZxg
uxllNMQ4WYviuGtjglMs8EU3It1VQtil7LPiRUv0QLYXuuYR8xq4+zx6uybJ5Umf
zpxfR+EsuUfJDh2VAckfVVx3hiz62yT8PUYoSbBA1RY8MqTPkcW7IygPAP6XhW7v
oMfeZcc3XkJro77ozxy2/xYK3URerMTWuK95/EqcViCFAQeQdMFnx/sWfAs/ZkCO
JeMHY+gvxMHuo4htNOyuXuXjPD3mgd/VWbV+K2tpdinVB25Fuo3Cmvumq6ENtL4p
O+jkwd77B82KFuu0h5q5UT+cDqo8BMfLSYU6BrNP4dPRnQrBu7LzX6BMXtbZvUaU
ghua0UpHiIF9SF6NMqelypzXzRZW0OETlOLd9770ytTWa3Az86iyy5WPYTF4u5fx
vzXwwGBgnlk4pSDvPq9Gsj6aOXq776EA9y+fUxwzSeGrQETaBbPE7PWEUqwG2kra
ZL2GMgMtIKulPFLhd/wem/O8YpFcKjVte9MM3yvnwIwKyaK+cXNA9be3In6AIk1u
5VX1HHk2JMhU29Uoe8tJV73w5ayR5Jws7DfUmovUe4gmQhdim59X2u0TKq7Bn43v
rviVnqUO3nLvfDDAs4Vv9SyeYpXGqqll97yEzztDqSQ5W0MIrnAdIfvGvuHgticc
VpTKWh52k6ZCu3DoLA7JZQYUftsGcEL9qYAKGuQV0bJmMG01/o4WG40F1w+vKQ6w
o18NSKuM+Ub+IdLr5qM3BmEUGrMy9/Eabr6x5dvBBbiPTXkJIO46vWnKgP8WsT3I
yukNXCAW+HBhpGgwGxyeVUShvtiD0GRqMjqajBqK5ikitUr/q7QtPvY2Rz7od3qV
GpSt1lqdC3YoDA5gsnw8zS+UwGGZNu6HvyjtqxMHqWG5sYxPxOObbA/z84HhDP4q
+U+Nxtls2hA7lU1gvQ/vOGj1PwbLV4UzDNGj5gfnM/FCJK60D0ekdFAO0H4ahWh3
Gre+8IcmaXsuxVzE/jFunPAoXmxvfGcp8kQXVqnRqVQkUXIt8KKJ1cIlhjBvEM/b
BY0vLhjyFH6gG3SdhIDroIL9v/as+FyE8WWGeQVS9ssqOzYRdzSWl+whuBW2iZYE
gEuAQF5uHQkXoWEP1sswjdznhwYnD+KNutmBOni/aW/mtnNw34hk5MdIbaSkw/R3
aeTQkr9v0aWre6DJCFgU7lBuKDR9ygGq/o+9hVUXT6KvcKZb+G/kZkeMkHu/THS3
cF8Oh8lcNgb98ZSHzUPcO5l6bUnHpgS9yCqr3MvV8upNjKCQWYT44MWhHsirvVSm
9+XP9qhnkoUu9gUUh/wHKz3dKqkwee0KXIuuV8ENfONuHn28LxA6BhC+w3QQxf1O
IzaPexRbjME6jzLbUGyjR2ZXoFjhvklKu/JxUyGI47uk6xYPAm3kM5gCcqilFsc2
a6NP7JpWrH2BOPaKWLCR+SlFgsxbxzLS634zU1NMMxewMZ5ectagbyirqTjZOgqK
te0SUt6O7+qTattqkAxEHpVEhYLf/WyonWjifPe2la5yEn1rITsOSG8TSHP4pvCN
WYAMazJ6I+pZgngUU/PNVd4gdo79vUxxEs+4puxC6hfoxD6q9YQN5CcOdoaL/+G6
xcmMgDpmtJ7kh2a6NX6FoH/TcEkbynzqnaz7VCsxmN2Z8FoPoK3aCh6h3pDVv3KM
2smtlj3WdreecB3fnNf2GsJDG5iiqL2TKnxxiEjgHloKQyQQeQU2C2qyib7dUoQH
xdtpQyLISiTwWnEqGv7e1HBhz07x6xmjiDaJK/XtAiRsqd8115wR5bBgg+FqlCCA
SeMBXEtCVmazDqZYs8JV3j9mWqWpv42BA8yYPHoUMWa4AhuWDg6G2qMMNlN1ISsP
kdG3KFwnYesJ6L+b7fX74DTbWU4qGmRNZVGzLBed3P9jxwM3d7R5KrDidjWm3SKV
MbLP+kNdlHyzE11hnLpOo9DyLZcgqSMrPEFnylKQV7Bne5VfHlCM9iYpdV8zK78O
PSFN1A6e00nvcj3AAgPQ/qTdT//1U2GZzIn3oTEbN9+QYZ+P0CHSDi3d4oFRIQEr
miJ+A05CsHGEUuHHM1Na6c1ELOuv/LkIrFnKAkZ+7uPzdyn4i0K1wQbkj6Kwtj+m
0cpts6BQ+DGkOa8T3MYRxKmdl5IBSzIu5bIQK9sDKsT/hhheKBH3UWw2u7y6zedC
6wiOSBnRKk8fWlL0i3k2bKlZo3Rt+TrFbv5M3oGdJZ0wETqmfR7P0whbNcnpw4sd
AX3eMeYhfozWJ4y/EUUDc1bExQbB7Zaj8T3ywlHb6TrZhbRTeEu+d1tVodc1Q38k
r3YnxNWR8ZTMP34QR8DRU65Dxfis/vr3eTTIzlT2EFf3bkDhqntnwyaG79jVnfaf
ETwh36+6dxR9iSIm7iayr7WNbj9/tGxdip/w3R/cmnvdgoxUa0DqsZbY/jVRPGQD
IP6zth1jLlcevlTf2N86UHMh0Lx5wNpI0GSnwwkSuSYDKaDmvzqkEk/XQrh+TIN8
6+OyGiI8Y/+coloi67YaKPd4iwKnpQ9zEIKDm/RDSy+lgsh2VuGk8cPA7g1Yngjl
nZK9k3m6i5zFRlENBXsH2sxSxzsPqL7hkj4Op4Yqunx2myrwQUKrfW4dPvgsfjOQ
j/1LPlXELWwmQdUhs/lU6Xi4Ug2MgrrEAnQ9gi8ain1MPFrmRcjJoy0vu0gqcqgZ
NTdB10kOxl0mTiBRewM88nvkGD14RrickpE6KnkUnEl9tZigRLFOM0+ye7o3skzT
Jb1sSSAQjxdXrBpmAi2RvMioJ1MyLK5AP/NmyxTn20WUprLncrK2Jh9QnQ2RisK9
5hgoZYFmjyd3HDzcqGVA29H5cbhVbkDU/PZCWHTZuL3qF/5QJchdnmWzJ8XsPJXF
7Izab3bM1Bk0WPm3XaZp7qcdDFgdVq4mI+n5clIWe6FVCaZEGqpTKqjStbxmBi57
mCzFYwLzrTN/KfeO/ZDZ/kO5y/Hq2gxmY+HwD9L8qXP3Kcbn064Iwrq1rayA3m/x
AkAxyFJZPXE7cdnxisJ0hUqI7bbVxWFOM/Dnc9RGYukHuCulnuasyJp15YULgtAc
D6eq1IXdyCdSTMKtM6Y7XekvczoJwqeB3LDhkB6Gp4su2V8BA3dk5PqPCwl/6V3G
EgienWrFcmVX/9dJECpPoFQd1UW0ZzFLCaQ6tOhfg75aVWg/F12s+FiocVMxv/Yq
2m9RKp0KCOfC7CPGI73fDRQ1TXoTvFIA02wAroDPakzg+9S5qhFrjwy7uTbGj1vR
8YooPMs/eGSLIQ+dT3fZcV/a5qOL7kEGm0+dAPNtE0PhIkYSzAVsPlvLjP7/K8CS
XSaf2pvVA7tgXSqWogeTcSdGG5aRU65r6jnVw/6Q9uutl87IJAeNnzcnSMzaKsuB
aH8+ue22tnfkfTIepHQhGnq/vRQr2dMd2tZ1Y6ZL3PPkZX/8o3RExQ5DUKPhXEaY
xqxfcREV+aYOJMTc7TrYmT3SI+YXYcj20jdelfFltxWlnAClvJ/8IVLhvpC55wpe
z4tk4Wbm5/+d//NVj0pHNvmggj1qZ5b1OcG+xQ5tsm4bS0ouM7OBYZas7JTYv262
Z9scqfDtNm5GjqBVfEkA4z8BqrujbI/uJAgnEZsLcSIXoJxPZPQhBf1C4gYI+UUh
3RPsqZlpdwZPlHg7pIel2OdXzoxNbfdc5lCnlgJS6IJV5Pwwr1SBijHNbOJwQUdf
N7uws3zxLmLJVsAC1UOIY+cxfM5mg5hR/hMCcU5NK/n5uD0/CIDygiEMF3r1ruHb
VjAK37jwv1xN9TWsZEuskoZcS5SNyvakwNM23oRRgnKADFHBU6huo1XONzD4vLkY
KUO7h2xrDSsuEHHS9r6xAwP/wbPYVmPiEdDw3Sp1SDG4wHldOn3ls3kDo2FTCmXU
RcGVJxZfSpffO+o97hGrKcPAUO7VzOGGK0vvXJ2Tt9Z0Vb8dKuti4v0gIs87Z7nm
m4Xgikguar/hTEHgFDtdvr85yhhx7iyLgRH2/oJFaGId1lnxJI3YAIxIz66ArZW6
XyFE5NFD9ZfE2HXfsmpTLYDeFjhqiLjJ5F8DPl6WXIF8jvNu9f9Dep0nyVu+++p9
HGCCTVfpGdaxx7ySUVn9tGUrMbAhu2TtUxdqpPaleaVmpgQ2GxI78eXKlSYQ7+lL
3SyxFvhAn1iHxDE4swjahlkRE8uFpQiS4SQ8oREbhWJLX5//CGorv2Jo16St8BDk
9k0bKRT6xc/LhExVaRv91oezxg8OejDGoIbupyTFLlYnST58FkzxAPoCBbDS6x8r
hjtBIixf2qX9c44/DFl3/DM3RW6EIibU7sDWnGX76BwXsZ7ljUWawuPT+sMvf8bV
C+YUbZdgGwWRJKYb6Xli2NepokMJfMPymhTg0TaH4F9DZfWo8oxijaZMllfT3ugi
54WNHw7v272ed1XMom3cJSskUdNMqvsvnYa2VAoU73+1QJt25cSxA5C5XDPWXZlQ
B8aP6H8SCVGf8sXBZd6DT86yI8o+cjjEIpgUXa7Z1Mv4YNzreUelZgsVqD50HSNk
kSHoWCTFgWh1FqdNMdV8irCq6983/HHKtVqlRw/cpODskqpDKcXntwS6lt+x+Q/S
LtwzHnMFodqAu4g6l2QmVJ9Dh1mp4lF4p97tYCzOMsGklE8wk0jBiuWB0E/Zg+TM
dFd7aa39cNLxeYUOWj2iAXmysrNmAfpwDD+1jhyaIsCGOjVpZJVcZ35w9y+2Psi1
2PKJUcAXEFthxtKKuo4Mc507/dSxT73xjOGxCJsjwuIEvAWdRA7OtMYbdWM/7rv2
8oBrJmi5cXZ6s5fROGrGyCFBH01Ky4Lri+q84KntFmJ3mFIyWXUzT4oSCs6JVgYE
zIYN3m0lnjHj4YE9Q+OB8eJnOO9CjvNQSfNloqPhCwQKTrthHkX9UgtpLFCF0ZyF
H8x+rXQPkJem9PTjMqcsXeslA3fVOB4byN0KmxnhabEOVHwwliiuMJo3aRfTk8pA
Oh4wVZ3BdBhs2jTCyDCUw8vvKUnpCJUDoNKO/VKnZjmSfkj1ly86Wd0ssZaem0uy
ws/j6/aClr0yhxvGg2MwMA89qHGb35Ygiuxdai4lLo0J05is1zVaYDrJ9Rq8JQNt
lJqyxh6IEfsSXHHQDhAVJQZN458a5UaNxtjUuyuJP800dMX5D8+YE37xszmCGHQt
zf1sucsWzxXlFj2EUqB8I/oeK3FXEvBL+ijVsLdTfZR7bpgCF2yFBFKt6TBKq2VT
WnnsGYkVZtShsHXgE0C4Ny0W1qDUd7S1Hte2mQ0RucUvKs8BfwKvYZ2YYBku4F7q
PjHyijczM/SNQEckLGmjD6fOzZzAGct74/AdRaoiJ9dBG2RL4xvXmI8tRbph7RkU
DXz6C4Q9ZznpQtfjI0FbEuZXnGkTJrTs7vKiPVTGNU666LEegYzSVimlWjSu5Tm8
5XZitFsZpuCpYjibFFrxEE22QccWcAye/6fZtrZ9RZEn3GvZzu+dUHHE7fV0elWk
dRcJjnSS8AGeld5Wi8Ec7PzReWugMkoYrPs4q3B5eWbzUWeWSH4fPtBodEyRWe5e
Wf1ly5w1hw/w+Q7aeJyL9I2Q8uU0awbcXDemVUGgRhh5GepM6TwY/wttVoSfJ+Er
LKMClgB1qhshqqnsY4CPkWrh8oZlsiwDb2tnwixosMaYzV59oBZnRzUEb8RuFaYl
4apHNfGpDZARHP6dW4SgRMTHRVy1lElm1B8jm7CUOaHhMmcD4WMlsu/89ASQ7kVK
v30kenAWBov7djusgd8bj/CkPQziJ8KG9a77sLRLcUGDcuLOO1qHus5vjm3i7hEw
idETJcwX46ejKjC1wdjuoaZmELqnSKmAFgPLc2xrp7JY5Cav5EaDQs+eDPBl7gx+
rkqARtJlBvYev2pD1gEMKpmZYIkrnfmwPRxqoN2WdTTcsWmuit4FVhM8xW5+SQLL
jEhmX5wIO1OR59E2qr+hQriiG4rol7tdRi+TZ7/rjVNMIDZCbLzbIGjmlBpqwHmQ
1XnVVTXWXaKfNyKtmH6dUuK1Z4G+aTOmElvduMJvQTk0rt6Jn3M0739vl64cSSDn
H+mSB8JmkeYbuN0RbXqtuDh9i28Jdbgi/m4Ke5T1iFVzzpI0HX3fO9yOPurG5/jl
jWW/4Tl/Z2Qra78yByrBR7A6gcE1HsahMthsl2H/BRKChoFOOQ2nzf7a31FwsPxl
9KQBTTp/Q12WgkdIim53dgZRXzcvGHMPMPEcbO6EaeF+e8dB1Sf/GKQdaIbKdvur
ya5/fcCrZPK1r4wit9EAnG7LHqlnKj7qg7GzoNfvuRGa+fmQZ/uPYgbAnX9qwtcR
mG6cN0hsrks+K+58es25mzso4GsOD7+jgiJU6qANEfh3TK+Q34/epVqWYU078L7g
e4h+DV8082x4ebT2bGWc2fOnACwVmADRsOyB2AiH63S1bMRpMbs1wKqzx6P5NJj1
Nj1LxC+NXd8PYrclw3Ez4kYA4bKD3jyzORvw/qcu7sypaFSQlBR365loz5awVqjb
hSX2J4F4qOrSz36JPD/7/8g4m7wvSGrF/FMrrW5/udgMU4aopO9iKIwObJVOz5Oy
lD12mpkWot69TX4S6h/xK+IzpvhMamfQXPZhlayFsB9iiSP2Yx4x5e6kvaxt3cnU
Dc3/IJstgITQ5vuUc9+bnnEp+FcSZsXTyme4TLQvt2EisSgsjbtVuusU4LJ9agAI
/d6kAjqThjttkCDAEV+LSXukiKzV7TU4BF+d2X45/AcrLXnrXHA5J9zCOufC5/VQ
LIG/ZFeusDaKM+1/T6mTHKzqAj+UiPYIiPyQsQzCMT/XkXrRppYFZfCSJ4/SWSdG
vld/837IEcjLGM7Dt0uFNLBYQ/Yrp4pMcr92h6XfjSUJwLdoZ/aS/OfTBgEFNWkC
QmLMzlJNt/g2xrAXY7Cv1Lfzi24jYJrjvcTGlGZ6yGy7PAGLAWo0f/GQKcQDiIau
XEsaDbK86THyOa68xLAIfxYoyVu31ofCELswii0/a3jrdeLuaDgiGCtacTFFGvxx
AHSL4WBYZ+CxyrYEOxoprctR6j7iFu3TdUwX15o5vPvckx60u4Ai3Fw97LEuCKW0
J5sOgKj42f3CgjiByyvdMCu4m4esP6tFkPlKHXtxlGAA3IsvXRlsEEaKQmJ7N+Ws
QgNafbT7QeD82qEuDN0SePQunhuRweUdohfaYc0JyJvHA5DCOtSLdZsH8Wu0LCYJ
zzmb01ej5x/zbo2Hqmy23GjQ7Pr993Rp/+84UhQFlvAcUILdPZXNvHPp+4VUBFWy
uxtULn7YlC8uTFAg8gaUGM3xkcab+l1A5f6aFguYRcFoVAnX+3eDQZk0CdM9v2Jh
uIjQa09wghGbnwXEgGenvYIVZp5DF5KYMi4t4bv8hymUWPvPUU1zKzuusn4gMYY5
BesMFpanw1JJWzZZ+tLEYsJKlrZNwBYZmMUDbr4B3c8ZC5E7620Z00Byqqxkp3cm
MrnB39Tq0AThfkn9QEOa9Dj0mK+fgua/354ddFIBZoOxa1CVNgXRinefZCg6yrI1
x+5hlL7sJZVDrtih1iKsAFraDaQ1B8uX5b6DjJ9Q7IlbBNQIGdcXZ+SBrwLu3/OS
jqp69/d28EdMCiwQUapkEmM4elB8mglCEfxft0Y+y6A74eQb8DCjWvgw4HGh4CUJ
ytGMsd/VTPzQnECbpJYq0cWLisD0QlhjPPYQIPEJiCi9rzyI5/3mNWHeA4MBtlxe
Pz5pePT1oLSMWLqFdy+o1e0ICE5M14vLuFT0g/6wzj2hZmOhBCRRcaHZCNgAuIC6
2z63K0k16yWZTCfq+592cEM0Pq1GIiyrh1Td2boGlhxMcmPcr/d3y6aduqTJZMw8
2AO3qBTq6LuN9dIMNKl0ysICRTAIHbOSWnx7bNsCTxAYZTsbUel1Jjbh4RFjkW53
RmH6f3Vfpw1N7Cd/mIyiCjsLioYyuwfEendYjFmiHKMGj9uTYGndfwQbpFIPnk5j
h53WlNj9RsaffQuBjN1CTTJUmciVZP5Jy1RuHesRNcViBfZXnbMFZnrQMR9RKo/f
aC66VRKJlVb6Awlf4vBt7nW8ql7Ky11SIlr92S3b73o5sixbI1wkk/dZITfPbUiV
ixKofKq+M/qeMxKqm+qeiUEvzwQjIbaaK9fu0CZ8W1iCBf8YsEcqY00YcYlPOD5c
Cnp7vGJXQd6ypeR3BUrCmhbO1aBElvTLhwWgwp3BQmEMUbRU2XRzgDhkae9k35P5
Z4KTnYfDiphbBTK+O0P8memrr78OtJL6hbABTGsF7aQ+by/aPG3CFTA89zB0ut+K
scLbH67FyccfM6Ye39CfzggrUuYetCdHxxWSQC8NTZ6j1Mt+3fC8LKLWwiigM7q5
u+J0qMbP1BEgwmDoHlG3xXXoxYuUUda/V/Nv+7GYzeqtaU9KnNA0/KdR1WEHw06o
UYZGnTWqRVk3GmRSe3d29bkr+fGCJFBsEyNHlQu+bt7taxUH8QgEfx6k4JjIFof/
gqR642OLY1kNFiraa2bMyQLtT8vq6AdIEi3j6H//otP5aOehM924fVG6iLYV+Db8
/bAgVQRnSx7caPg/Ho408cvQxp0KYENWR8eDEeDCCA6L8oNWIp8lgm/3yrIrtN3+
XGq9vqD+GjTEifvBikxpYT6fa/Yut1h212Cu4TQyZ8aEeMamKLCa+Em5vSkGX2fH
URLN77okBacuDiFzh3EGEGQoUM5zFadgWDNAHWfvEUNcHLnFW/JGgE+3WRRmTFj9
vyJn4gi/howwo85/iwYL93hqZlRT1Rfs9yspCeKYEGSyU+JT5DpyVQmDAma0RmJJ
0FJAiOriMHg6JLLpdlvGWtuhp3//HtcVBPAZqKD5Y1P3LnZJRkGyxuawdpTr9+HM
q6/4ZhYxRYbUhUkf6yQO7ZhqNpoglRVb0yDEx6c41yDcT6Ug0J7XKwtGs4LJJEZj
ZvQCBsMBHgqe7rQWMB5nHV0ruBVlKhoEa65Z2VWq4F/7DpTCiW9bNIZxg+TQiBP7
hxyaqk81sIQVd5oOb/Y93iQ5vbNTe4cOK8TK2Q63gKMWUh2DK5tt3adj3b3q6yQe
CZgMB0RuAGkK+mouGePf5pPsu3hObDZKxHvz8M6Gad5N0Saktth0Sba0nSftlKz+
NcezBLk3m9uMCTfBGPdyengVzasb8JDUnd63joPyPxgw1j6eEwvpQqdqOURDF9dB
TXVh6kJIcY692BZGv1JAFYkkzzL6lFfeJyXVEvzjhZ7BQSQqzmjqcBODBVNlxUSk
RGXQxwrUYwmA6SuXFAZGrUrNYetu5XeeOMtIYieBB4E90i0U/0RISvl1VB8wFTsF
S6scgg86onQHxc3liOp7CFrIhqtB8A5w8vCU3g9ttNF0jaKoo6Zg6tXPdE3uM7lQ
EKmXr+SBj7hkpiFoLV3q86I8V27/k7GsxSpZtvIgkhb1FkXMzEj0aNNgXc3W+PIw
eWFZarjZ/nZjApQtKnCSy8orPS2mrqh9E99fo7WcctI34ktMWC/NZQG5wfuk6ehB
5Xco790vsA080V7gYbkByQ8rAbwPwvzw/fUoma84YMEC36vFgqmXTyhQE7IX3M3Q
ShAYp89LAVaFLsG+krHWSkLXWurH2ZbAexn6XabFIfJ4Juy2c6CsbX8qCRjh7nWb
9+13hreSpGcKHX56Y6VjPEUmhxN1Sa+9YbWfU0nZCX9peSpSM6hrNZqlT3glMsRh
YEfe14n+IlvDMZQodsgBYSPJEDG3m8j1W93FquG1Fo4r70c1JOovPtZmUS0CvP+a
KA8UTxSi8evwJVdDwbDZreBpPHkPsb0DPy1UWlyz/Kj3HS/itsRcsaB4J7ojP6FG
4mSBQcWKytbJ9Aq+UgoPiNKS2eolNT1uT0fRRIIQFz+A1oba/ZbvqLhOx4Xh8+UR
iyEgKoFz2ZEz4R91M2xEzak6b3oADIIGe1hIdP7N12O95vx5vNfJOsdoq012KXC1
jDkK209M+YKImfKtIREs02UQdtB8ngy1Z0xcWWU2eobMXHLiYVsxbqBypGpfBuOc
Q7QOAsUoCKxBz+toeKMADNhT/950MoEa+J/PM6zvCfc8sMTSEpBkXkTrOSXFFzBb
iUF4wZRu7645DsvdIgWID0liKDgVrOFvsAS0O8XxwJhWurcUyaCfjKH9EYHz21nx
R58QTsjMSLpQul5dwHd4gZF6UVoKdvWFajfvBiLsXSJv0UE/WTaufH3rVEiptFJk
ijr+BPiRz3qa+/1Z55/m2cQbrHEVJmlOx88ZisEjNukCW5K828lLVUCgG4+r8AIP
zyo7/Zyrf0jNBuPNpuA4qfHnAGt8d/1zvSmzpuJRdUC+i5LpbgLnDZwX2kJMwc3S
j5U27yDwG3JylW9b+sWt8ifIAlZkVSxQ2KLHosXkNyCKLtLalHj1mHBDeshJjcw5
DqMdD9eDimVvIGntw4nGFAS1+qX6JxkdytqgQ7tR/yySpyM5oGqtXAA3nTaQsIPp
mv8UGvGhwmrXLyTQ0XM5wrlWPeGb2ZkkNzc3JlrKPTQ/Gt8v7G0F88OOtNho7CEs
04PS62KQRyRWzFPWwL3ks5e/XSS4JxDidCu+eQi62UhheRDU17mIXyjvw00HhwR2
M5K6mP2SyZblI2n+t77z1UdTkvNwyDBfhgLtxawPwMRuPb6UkMGSXo8vR8YxYitk
3khj3qbPkWF2y8APnA2D6t6HFYYlMGOgs0LPRuDhwJMUktG3DGLqTbgfbFgWdrhR
bDn9laCT83sn88q+xSDBxwWcs8cHII3zG3D5lK3Yl+KEdDa0g8/Pi7NlmK3nXY4J
qb5eiPAvPrOPmei1GW6ICyQ5k5+dlhmoZeNtOSsCahpFyGCCM7U0Gzh2Ib67zM9V
ptN2GGKExMZMb7OPV6o5LcNG4Uc/OdQRYt4gHK/pD61ddd5N3Lg7/MN8wmt+tkhN
T4/whQ+Qc8YodsG+oFeOEuEGBuhWlgfFMZMGLntLWUEoFWPRMxHlK5Q0gxiNojo6
2d2TNCcxehgc99j9I9Zr2s4vPeboYWWJglKVq++ZFS8Eh8KXY6cy4+sO0+DlhezW
AYuBzGdoukovB6hOUWyGo85hk0qJ5DHu5yJK7Pj9CbuXWs6Rc5UYnNQG6MBASxKY
Spwil0Tju9D2CEx5ka7N19RAexteqhy8YGCtS3awzC1WHfJXuwf7u5x3nzITX+qh
ke9nwNUSGhNfinRr+VWBgiSXH1Fc0WmNAjVGLVny1Hd/ngPuJ/1+B0iuwzPUKwX2
cSKiIigVUOPtL+K/FpXW1dNWmRdt3Z4EAnvtHtnNQIPmQWdLag2Ofa7LA6BawLvv
qa8V0qBvZSXrYBHSy93JkLelcnCx8MyUY94+fYVIG8us1YxGFmMxEe/MOMRKXHKx
MzXhcJ2zw1ZrYYzaOOt+FkKDz2g2TR0T2XV8tqoU6XgdTgJhwINTFxMIRjKRlBPM
/SgkFgqYuwPD0uyjouqUiTfqeU/EFk1jkZFdZkcCtzoIWYea5IXXVo6IYK2IKhV6
WqsxTGFb9btMIFUHUFxu2YS4VeP8DQlPFR01yb/9OGZhKfJEAV6dfj1cbR13phSs
66woSgVIAozSee0WnuQYvOb+KXh6ECKZ2b7a13Y37K8ap4xtHIFJcNi4DcFeYE8L
e+bx44uH53ddHuopk3sv0nBBX2mPU/FYB/yabGgMhlC1FNxz1U0jlC0HPJYHjVNH
V0y1Ml5pB7fxef3+aMsQ9pVA6wi//OTGh8kJKx1oWkd3Sz6YVqrq4ThAtUdH0bKU
/gmwHNJMEX8N1b/2TR+OARpZ+8yjnhYIwF0nszxxKcAB09aztQqIbbJVG4B5Mda5
qorXnITBHivLYJN0N58hVzmsh15Y8rTG64EbcQcy4cIJBLtToycUFL7A1VGJQ04A
SKDpuMqnd9Gbl6p81hczDPcIk6L9W9hmM5jD4YcKjhIYz3VcP+J3zlydU4f+gKl6
oUNdofEJYAas/4cGdJaQU+2rvvH/Kr2zN7b3+Y6P14qupQ7iw91l9g4melPrhaPI
jMaxneunsKxncvagtWPSQKqvHoHSI1SWLi9NGB3AlGwhDfoK1I9SxbM4DcSW9JXd
ezq64evFOvz/+lLlmbgBbuoJVzB6ApS+sev1RyVvNywo7G2IdK0oLHw1fnvSVlqf
sJC72ID1omKz93RefizlPHiCs0y48qv47n+5rxxMpjejVvcQkzMlUFn+FC6FKNW8
/kyyJXxw7cmBCgHybtWJjzwS6sMQpfkLr2BnsScqT+QLWTuDHNwm0N28Bbr+sb09
rIZ8FmHnyWxh1roUzEECP4qqkaaLUP+4rNSlOURbYoOE1zU8+s9uPGKlYKywiFdS
mrd1cBVxT/bGdZ405M5K7VQ+MVII9a200HlaI8aBtjycnJ+bNN+IzkZv9MRSt3Yh
ykDDyxvjmvYIp3P+754mdkvoGjZEdGTBiH3m26eTwOYC1rIgBaPi9dH1pI0WXr2j
cOdPAMw1vnhPwA5Ifk0L+Iw96UjabVa80tDFh41RA8DObn6JhwxJi7eG+p+DTbGg
65FQNIlnWDhHZ3AJ3zCBf1URNzO9sNIYSWHqPnRIOuqfnHz96sqJIGrA3kn5fRea
Mki0O/uQCUEceTvxsGp3sBY4dWSRJ6KiQl1vjvr6iaM724v1geVdJHSflhbmrq+4
XE6Gr0Y5bq1K8e3wf8qTl0TfuWrPflf4jwK1fsTFsj2vQ57aMwcUk5jR9moSaO8O
NR8jKlovqzT95BsE7a2u7exZX2ynOxCEMi9awQb1z3VSLTugoDJ4pQSYuKLgPDew
VPKthvhYpEsG8J+/0RL7YbX09PvrMucC+xCxX0fxMp8ziDnKGhzK+DmdALpc08+2
2+EjaSHWEacJbNecUW04IsUEA9ywiUk9z+6BFr+CM6RrJY4xSNh4CCAy+xfqhezy
0NgKyQCw8fCZJFENaInZ1CAfxNgl2PnekP1G3Fd33Z6Q2m9XhR1ar+HsuyaDs5Jh
0Hdn+nfegZOsGPmaLOTxXZ3wlnpjvbvFNYti+JFoQDsH0MTCwP7El8Nx203XEes/
Y6Ao9HvqKgKdNuSNNed0d1SHzEKoa906leiyMdzuoq5kvwH+4RRemEs3FYGnWs/g
+i+5z3+oDqYxtp3vygDAu47B3yRgrNC6fZzcpa2kTDxHhKVV/XIWMbaXHKM/1PvJ
sTBeKThBDYWmqiWjYqglNXdE0PpJMWlhxVonpeJYmjlZ/KUWhJOvXwiylgGWU2aS
8QwKj0fOw+jrZwdh/DXtDfQQ2FfNKQnqIxbN2R9O11hRTAAk06H2dWeT0kbfWnH9
Af4Zx9KSbjxQ641Kb+8Ern3N8X3KZVFFCLY3N3sDjHPWvg6Xow/HNj1TFTuZqz7I
tyRaTS76b3V3nKjYk1E+hKZ339wwr5JindYAowGVmA4UMiq4lHpE7K4DY/9C2olZ
SZzsoGuhhfoqQiOPQVLbHwMEHAd/NqV3+On1Eum003Zrq7tLRxmsEQczuYqYx+Y2
XhRktUq+I+32fGXzgKZ5nWPpTUcJkGt4ExEcqo1/0yYXA1CbOMDE0HLt+CD2ochC
EupifR4/kdCMHeHEocMIpjFfMF8W3aqCsLdHVvYptft/OhIbrsim/KUt7CDrvVbD
/RsWXwLDQzJHhcVWru8Z73B/5e3cxNg0sdQTE2BAdePiX27/IkOTyraeTq/U5ld3
nXsFbt3xhxfJs+Ui7kdrsfVNgXEdTONsTZn1Dq7/Qz/0QP19sC7pnOdOJf+uhxzv
6P02Ec+8bnSiCUwXAQQ4TYrZZsU9b6n7yV9aEYhm5/Euea6KqewlHITQAkXi0T3q
n2kek48kARqTOsaCxXC/824BTndnf+dHcVk+DUR0U0HEujF4itY7RyvuVottvsmF
lIhZj0yxIL1MKu2VEZvouPOu6TxrDPenGWRP3MEOZFqpA+1l6Xlv/pkyBKu12zQr
599VgUTVkd+6xsqTR/eYNPHaI7OdEvlusp02PgsxPmMeeu+C1J9N1gI4j/xWuUqq
tG03gFXXBV3oHu8mh9sGnZg36/WMPR7dU9GKM/t0TIL4c8vDWC5EG+MrTb6KAGKH
cc9i9zU+A4o7R4CYLi3IilHodXMjqGJ//pPsAhs86OPM3fSkvEkbGKTQi9m0+q+H
A7xTaanR64pj8MXPxJrldLZyjfq5kSxF3cDGrQwLhktfu+cO2rkqSrzQy+MqHPoK
8f6+qdXb5FioWw2g2eT0uqRqdmQ+x2Wo4tDawROyXoX8nGJsM3WR0HJ1kBAkpS6T
dg01Y2xDGfuSv7/idSaeCc77u1LEoTeMvCJLGllIG+K4p34JwI8T3q2TnZEQk4S3
ApORoPssyMPgPnimF0BOfrJXO/qJDdbfWf8HteIa1Z2Ot23R534b3gMkVifJpfin
lnqg/boskPQKwVJ1cpU6WAYG9dhn3rX/eXtBFXUvAujENz5TRMJjfjQLER/N2mTC
6CNYtifUg7VsRoR11hBUkhgRkFDhdkms24r81jfB8zhcej5F8MebXArffXBWnkBX
/pjwptlk5PDYzzNi2YuTKzlxXOyYdeQYZg7SY481kQfTQuMp4UOxoXPlHFLiwJCm
FEAvlHP15yLO15ZE8PeCgtDskgih84wHOIAfftNo50k/sxkzgHqeheZT8Cfz+mzd
5Jpid9cb6UnOfniazUNFCL7RCXhfdQF8AT6yil4vHtwaNfaLMg3mgukld6QMlnNI
oWGuHkWjC7BsxK8bNql5bPvCF3Ecv+hGX6bQHdKrkSUUIgua8nbp29vUeoDmuzxe
nNcgfOfzkdzUkasBbFwNALAngKZjlvPaEqnHSrS5ArUigO//f8T9V+Xp521GtXMu
kpbHYN0PQYm2tmDX+UAyHvCM98qKpuKQDdnnhqDjKlPP3bFh3pQ49pRC1wLERt81
+qp+Ip2smIFrCDolZHL00sSnFezIVJ7slDhCwGrZPcf60VOJ96d8uOR2Zm9Ad4hC
U2Zlf07HGQFfxbhUqociqJh1ilOn8StOA+2jfjKRR4PAOypztFK44srKu+Fm2+B7
kh4BWROpAFnFd3pReajLJJMfc7XS2d8k37E3tiSBNfvCQY01i11hQ/C8uml9t0cs
odKeSKDB0YCZUWkErQaj13QVmEy+h4CBlzXfggLHk9JsOUZHM5YHJfoSMwChVtU3
YHHbMYnDBvr7RzS6gycgtGZ9aHNKXCJHGKYtob5DB00DYmF+2h2VHdKdFEEDWR2i
cXqJK7Cg5h6FLzVN3syQ13nCuhZgmN5jJuloNwshn3BUkSrLnKrjgLr9hHzaYD55
+B4R9OqnlgQSuuIUcmx+Airfp0//lChusZfNSmxwUYE8AhRtb1jlOHpobssaH72O
fnOYBynzbN3UeRPsGfFEn29PQbUCXfoUJ5VNjPJb91SJgNftSvfQTszAiSe7eOp+
kIF6yVbL3js3/MUO/WiaNbEmhRUj27vgvpA/k4sMGmcSH+GMGHCRlcbjYns/cqTC
8/aFfg7wX7U4EEh2EXgA/jYGCnmRNJvzz4Ak+q7kp4Mh70aEpxVAjQ8ymdhkEhaH
xKCUDhrg88FyX6RwaCNp1vauZb378j73w1LNM249zAxyTZVbTzi3yOLucL6CMYPU
FMsNi0vlvVK7ov01v5ONfJwzIB6JnDGhwOxEXDGap82iLerFcSNZr0Xv9+DGw9bO
mX2yQMC4n2ePP4L0QuBM1IhgzTzy4eEHNwSNb9u+cVypXQcv39KtX07qUlFk4ebt
ysemtfFjyOp5hEOW+HfNeu9vyCo68cjvMBK4JFNZxkhZje1/sQwV91yryXXmKbkZ
UCT/pNBB60gDqUwz1A7nLeUdFt489SnTZtDSY98iuMNGxlxna1mGdV6vv9tdwnux
NJXsEAhbdRRvhg2fG/qqR8gh3HHTuN7Gb4TVFQ84NUOhtLxALe66Dmcsk8XPsMHD
k4w5btuZzfkCxehvrWdko4pyH2vIc/ZIBYjQGpmZwKJJ+PgnEfuytEbw8nV4XYlJ
bh/LQvOx3jbgrwVzti2gMPgzWXBlvM+5E7UZLi5g9WDzMOFGu6a2CImD/6tqJI+n
ytaJ3lcmvrZDVlNlxPt8e+ReY2qvJ00txiV/3KS/ng0RsPuY7fb0vUkpIBwTNjYT
TOzJia02eRzKbiO7Q+8SApS1uuJ96iZt2X5ok5x/cM2POV7yKubQQmrKPG+eG3KX
N6AzrBZQRFscrxKliuvKxpUlGkE9yVH7+eup6qcHUMFBQDeDHpsd9fMbjWkz0hOA
HpVQGnCQ7WqlvbFJnW1snJzFTfN72bEJ+Ha2LZNsq7r+3+hePuRExYOD0JSxRmaZ
oqVLuCgPefk2W7XeJM+wG8CfITNnnYsK9fWmgd5bDqOQXX8NjOMTdQOtKKJ3OxqI
z2Pn6ucgVlUqxcCAJ0hrnP86p9m7nPjy0l4uCqygTW1iwjHzMwqYuBTwoY/N0KMI
Yuj0oxEKsNRXmQ0b+xEGmwxvxLj9jXz778yNJfodWZkj0z4SEBh7D0SBPE0OiV6i
mYAeSWywHUMSXpQDVxMZfyYsNzIQ0VMDBMKDRBr/q26JAo0X9rR0f/5eGTQR2Erl
wdeqKpnQv5R8ZNJrzUElSQL4VyuQ8Rs43rg1xuV7Eafj2KSFqbXPcADSlTjEqoGh
cz37FTM0Gow8rO1TnAseZRLTtNcWleAGRYy2t4ELi+i/AOf+Cl1a10TTFW2l2ayD
tqTgpXNK3cVSvPZqbp1CiTPTLMiUmwgSzPhuzFFitBxU01vSsZrJOxXkXCOfoxNA
CUblZvOUreVd0G0sw+F912Y9zt/h/CoAgzKq+touk7Qgdyd4GKFnLorMSRWDAhzL
hl1/oDNjhEAsGorZWp15jTQWfSs+o49lFTZ+c2NrzOSGlvBuqfepH2FwiLcXKICD
W1+Zl9P3ZV3cwixDYs7K5FYbE2P/q3aEUzEgzI9UidVovHPksaJ0au7FvevXXBdr
Yp3IDXdwAez5OYFl/YEged9ew4lv9sjH3w3U+7I+qWgBe9DrMZkLOA0CS1BEZWB0
TpAenT0P/sFONWr3DWFFSHbYEiKpjMqRyxJf7n09VQ84+FjJ19A+zlFzRSzgB1jv
OVP10cf4IvstGoOxfb+Q3Yr7ETK4e5JlLQdLUbAeRd3oE96HkBcU0okoDdUD88Ld
izDJcmsaVJdP3MW7WuRQl2FXKbPG7X85PyjB1tIgHRajpZg4zeMe4ZG+kR5mfHj3
+GefjxCV2rjy2xlkoGBli6EvFlF7hpe58B8yKZcucowfRKxvG9sFtCDBLG+ClKsB
gubzjY/z/jf01n6U/qd7DX+k5YlWk8PDHrlGNTyQ5/DfdlKbCDHztm60M6VUPpZM
Zz5tKfOnhIUlr9en3wVgJphsCuc09glSRTOPbXUrZab64i812RLehgS9nX692p1/
l5kyDpVZhZK8+mN+WOp4JBYuMUeQiD5US94WC01ga0u44hIeLzzZVAvva/0+9hXF
h/MIhxauym8le2bGmz6Ug90vst/XT77pF9LI1rHeC1HeIRL14Q8l9eY6fiILx2Y7
b9tuJsIb4vr527ttFfY42GD+Ydc7LphSWNxv/+SKmoWTjXvupT/MrE9PS38HASvF
nYUth5E4D+aD3yA+9Ig1smgdr2/UM40vLCbGT6Ogg2dwvd73vvNUgxnKufSpKsGo
AwcxjGwt/fE/P8khAZhpfyKG9UT6W/HO3yYZhsC1TNb2Yw1QxvVI4JCvzgWSEFMY
LL/SzAwiGVoKNS2aPBSSdr32anADQJByuhYuTY8ySt4guGRU8qFPOPa16xL3P6uJ
GUOjbc+8bl62j4zp/z1y+H52E16VghCRFFas9ooW8YA0k6X7ezUtENPxxl1FB5Rz
uObkPRtV5e/5wmMOYfI+iAaE4NTgnyPYSpfPfeKzGKU0c+FKwULZXgMQxfik48ha
yPl7zPFV5ZHKXB2jBwdx7nxboZBLeEZT40BRJHvGik6/IDZG6VV+vbeKq7h/AQoR
l5WGdmAriyEAe1oAMSo3Iu8gipSBXu9I1Pp8BSp/RFOygF1hrXs/MUVvv2fVsZIo
fE9e3QVJ3CF7541+xBM8jNkqUXwQEpXQskkLCdtRBPsOAmZnBC8ziERv3Xt2CBOV
Fy5G4PzIlYp66NFjjFDc31XwYV1BbW7tfk+a8he6jWdptGPpa3/R5Gk9cNfGuVbJ
GFaGo8MD0nTuJU6fH67kzn9Wx6YjK2rxa2U5F+jXJNxRUDFdF6MRgCtwlwwIsoLv
XuQ0lm2CUNC+jzNg6c7NlGm4HdWr1Uhf2q2KmlwLk6FGJHCyLf5h4Szal4aJDnTD
YGN+y+ZS32WawoibvTOB7V1tgKy9scDOckD6ivk0NE0drXYWxnesC1749F7YowhD
f08KfySiFXQLIGINWz/P3odz9op/W+HfadAwj7wrvTLYyYAbZzULuuHWnVAgUqxE
OxDsqpctcHYGnZiK01iuvB0E29ArCiHO8IHIgKWsZ2FPIYi5hjW3WOlfcFmCDk/7
iQdsuKZox/OYyMMARPVGLd8VDkc4wUmkjR/JlVhSW2MAvIvIlVyapYgR4621gSSb
UtSocwbeoLcGd3FlFyRL7IvdcQKHrDXnHwYZmeLtol0zgpBMH+U6q/LGTfuMV6kd
AsVekXVcpnc5DMOkuov4NNIAxbXr78I5OP2X8J2BqiPQwMZQBsN9tTgC8d8Tp4XZ
EAUEeC3Eyu5sfcnEaXZv4r+q1npkE7lORGL/inG+trwSG53Vp5nEciiPzPC2DeI2
63Ienlvz21QG2UVEaG0rjc+qh1R3b6XIQbYcrxQW3atIdqoTX90sgWBO6efSaFdE
QwhN3JGMVh4J4b5crI/Ch34/nARL9J/85NbULQk07b9AdR35QjuCV9H3jHJipCmv
1/xCVQ0HxMtxkuMjbFToFGRhg4nqPwvWnIEYvXh0HBDqrUJQdOTmPPk+StcWbFpZ
n9ivlB7nnyET0ez4hL3dOqXPV1pGRyi09aQ35tF8HkSpayt+x5txJbyAaztpwNPt
yCsQrZVbXn9VkqVsZNY6gNEYWqcRirrDnqwV01xAO+SY1A+jYl0kzQGSvGItf4fe
gr970XHOcommGLA+XaHBdLmnghwSxnTBtB9yCHgB2Pc095Z6m7ZDh57r0Q76Gamf
N9JKkgfucsRAp1FsH0EykFw8Smi7a3t0Rnek0MMYmY78nHi6IXlGwFL/UeS6W4RD
uz+Ztr14R7BIbKm4z7GkoHCJl2sy/K7i0H+ZkIefRLP7Z4ag7y9B2n2uALkFWv61
vUnUKNiK9relsr3D/JW95vKA6QMHf6I6aUpir6VYSMX1+g6S+ZVO5K34Gpe/UWTI
88ilWPuxI3gQMiUyOgj3+ZAEO06gVQ1kvoy2kSn/jDamaxHdbQ5rLo2lhhE5lBp0
XbB6NVzfJo0l+AqtODuxkhrbFkw4E33U0KsmYBspimoqDHfzQ2r0YVDsfc8tyqjm
EtQn+iI5g7T8WiFj5hvevjgptKUuqN2AHLQOsPy+gLkZr4d1bkIGo1caJywcxm4b
qAuexA6QZoOOrBupcampX3B5tBvOoNLSW6kxWly5ZvJS55N4yRMeRifpboEC4eyT
a003esOriliITosta98OP0c4kIdTsbmNRLL49yb5OK5usBBn5q0wVPyUwA1NzXPZ
p2HNft0GRzynx7AQBBZGChV1pS0phm+ilTTScPSbtkNRZliNR1O6ZI/P463/7juT
TvfNpgZXIpCBO/RZ3V1plV0otD6FVoM7eTfrhc6xKaGAsIJvtV649V/fXj5RS7yZ
qDzd/GgA0bF7giBm20LZkMmYnuPt95iG0CAqN+nSu0ihODtYSvcXZU6BGw1KJhiv
IvBZFRRniXXLH17e9zdRRiTZZNNvVz+O/6vPIxxS1bjt0IEibfVyhf5Vk/nZhlek
NJKzhZrc3PJ0aLRrX38aYiEIC/WbHjx0kvxXtTX3TUdA/wWqDsn6YXQK7nL9IovU
/HVOuyb9wvlibK1Ohvydn/mkbE77iSg7LTVwPdhkMQ4dgSamBiM+91hnuxqrfyW6
PoHn3BBKKjADn0BVezQoKTK/PLXHqsUJ/xmdVb0R7W3cJt6q+hvfm0HVBP1H+QEL
ss/2TwtNUbsmsADsq99VPa3D2qLswjQmU6YuM8ogP3v9gHTXTvZjsZ0/WEV8jGRc
cdkAOSmuqvWl15vNK3GkWslTOXUi09kYxES/5h5XTzJrej1L95mStRQzyZqYWoKk
RMrDaHn6YecMxHgrdnScSQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RGCpZLwOi9Dav2RmZjLGuXiKUjbpvJMj+5LJSZYMER8JWDioFQ33vwbjzJSwi5Rm
nEhgb/G7Fu03boOob1xLFNt5L8JgPwRAQTvz6BaqJupxI+SFJpqKKxI/YjfGl9+Z
R3JiaYUOY9XySFmLWg6kyhiiAzDzy8G5Zc84XXK7neRro9lhACChVtlyyX9vUSxU
5rE+w7yE/leytQZRjC3HITdG/MWfKrQoOPDx5UvL5OAxQOMYfUbCt+i3a3RENKyb
zYIqo6ZZPKmXVQR4he8tElYNV+uQ8Kw3cfMWBJDw4XeDzp6astKeLk91F+EwzaIi
WQ/UmmZEjJ2b99hkIUUVLw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15664 )
`pragma protect data_block
PbxxxtOtr9QVKppCp9/qsd8kQbyZFW2Yf1R8DYtTFFpFYHlcP4HMwvZmmzYVJhNw
zUNYE6G/Ud9ddY6RH6S/Q3aIVr6n/pGlARLTS2DHxAPZwLIDwFxF5K/4QWpv2o2y
G2icAD5inxoM3+iqKyJYJQ3hBvb6LiZn05dc1sT23wZ6YP00nybgcKoqourcbf/4
NjLOV2ayDGg4o9od0kN0vKRnCzKqKJV+RK8HyCiuDp/yjofZMqaD6vI89jjP3X9x
5S0AfIxjeM8wLd7PTZmOWM5mEx45HVnu06l22Sdb+/WskDdwWK4/gcInsNbeLxZT
KaYLgnlLljz8qhPvTXf+cq/Yd1Q3OJ31o2HWL+fzK6LQg66nLTygolQhGd4zPagu
yyVdlG2RAL/bocCLZEv91W6/t4j8CC8kcbJCylTF/AYdVtMdV7rM+opT7LUo1aL1
xyzJcTYGku7eJj+mxrvPCOtVnb01U9zO/HanvA33Qo3oguB+varvPpiwQuf5/6yz
U+aOM3Qj5grs7pz+lYM+wUvOEqFPsNpCcaY/CQG+pzXhCPsBbepvEGNIEqCzUY33
rzbL7YQKZ25xLyGTJlaQ1+w0uoDDo3t5P4Df1cs3Kf65XCUrViuEcCX1zr3n9D3U
PD4EFJ2yt1kq++KlSXalfwmWmq3wC3Jr5ItqfKZv7pfpIB5NMygHcV9WLVcNWF9J
3/ri5KtQ8f5qHTG7sEMq1tRxWF/JnXmiCNbAUp/JOhgYATLO4wTUi0pdLnpJIsYS
qc2yDKE9WvgUxz9hpUt9TlTflb/hUSa3mwsiWXuRjN47k7GaxuaBTloNG90wVYN8
Fau53N9nly90mwWSiuY4aiQJ+PZ3JVYflKYSoi3NRFdlWipLCdCgtzynZj7Xbx2n
eh6AvT/122ykNf7Q3zsRmdaesuCWSUciqI/lRL0ZA+oT9SpAGphkJbEXhQo4dcKn
317cT8eI+1+xcDZVQDk+XTaIVjJdr+d67X41R0DQoGnUq5PJJVtjc54vmgg+QLzb
WX6WTwMYQWLaXbyT6scxjv7oB805X4N3R2wreIe6nwTnO6eyzkNzwvDZhN0G8LAY
guX36eqvJ0aqHtZVe/4fnwgPYMy/y9oHgoeID/isariFSayDjT4gu2riTiSq3TPI
jBXI5iB5Q1q5LG3Dl/GrFxWPWBORRtD4Hw4gSTL4cJJXR07GlDeQ9L0YqxKrpA5w
Ew/SUXb1q4jKnDKCDLm+N84oB7Bs9jnqnIQBMWVZs7x06ZPz9DMaCltx9AlsRSIH
3YNdmpc+gGQYWAwk77059ihQJfJqBU6mVmqK0m0xKA/Bg6BFO2FJGkgD5b08FFXG
zADrcuOQucDOfwZr8XZ30oz5+ddyaZxoNgjOhEo/QJJwc8HfrWPjDwjDDDQJWCwo
P+jf2Sr2haAeuG7y1bcRws5bzHsgbxmBAtPpntPU5a1jKR+0GEXONTYQVZU0kMLv
2vu5YiPK5uV5F1x0h786jivA3NYAYdyZ/ulnPf3cyW2bUoF954+ZyO71MqtayClF
vAC1hBxEnNcpcWuwfNPZ+8hTtFDeVqP8n22pqe809kLJXLf128XDNc0tVMXyMcs7
fJzin2RAn8J7uY34qzcQ5scRxFOWJ7QcJbieVaAhunLtBEU9ABTuHR9SPrBwsfUa
GO7ztKCptE9sdKeN4AMB0jrLehVVmPi1lGsE05tJ8cHEBcVKdqJCh4duXzB43wos
jJxERKFtdGeLw0icecsokG0q4Fh2Na/G6HCV43s8JAImIH90/3NiNJCMj2PxhNvR
mTD6u4CG/lUEBk4avG6bTtCghGFikhTYBJjj/U2WdkUStti19+qYhamWq9LpR+I6
4ncv8PE3Trr9OfkPLC0uqLgPKmzRR6Vr9F229ERff95HofiVhVDvEgNvGY/K4ium
Nc7hxk+aBB2i9wMwAaXip7gsbIW5Og4jMM4kabJV8xC5tIO1AE+YXumSTXlSv7Ru
T+2FL/VViHZSq93MlrW7W+gMSXfBOifSvezla3TK4MhisrKihSQDM4nRC9rixgEe
8d9YVGmP8E2r30nW8SA6lH/JYHV4zrMULBTOjylaMrAkuid0WsS/nzCXlcIr9lMm
TVkPwz1R2jdoFK2FQvC6cbgyADBKhS/3CPrLoD8qm9KUsQASHbFj0WViacEv8Lkl
LwNjeqPdQR8oBp0XGnPqpyb9xpA++avLGRC9dYmL43i3e4nMtwsyJe8TEEFjEgfn
cHRiqOa3a+/oJ27DTBYg7rCiMpYB9oTorKIdlpQhWur+K0urhee39ffP+t18qVeq
V+1sMwj+KKJnH9cxzTzwET8JD+ILvnxeB9lhRW7v0MwJeHoA0zsX0Ukq2+p+so2K
ONImt9ttQMMWJNG7tZaoO2V5C61kR4ig8H4QJHraaqh7FKzI0jfKoeZK019GZ0Px
VvvnqPzbi2xI+4YOd5qIb6xqEBsxZRYg/EWkmhrIaNxE+C4ji73oYaj+7UnQ+kFz
R3ClA4FULNYgt3J2Yb2CRj5Dl2FmzcddiX7+yhq2owD82Lqb0Q/0ECoVuISGk7lX
ppBJvUggAKGEMKo51hCNHxqFq4c2JMjcfng8y73xGblvjOOgQtorKMlRnPm5nggP
vpDT1Li7RDymGtE1ehFmLZApgZ5R6jux7OF/k+1tity6ARzsPGi7MvIUzLD/XKZP
HSBG4c022LPpLdaVvxcJSx84FiSFjYj8GrvfQpJ6WNbJPUWDMsJYodCgYzEH0nDj
UzzJYK3Q3eLGvA823Iq1MAX5AJqVP9mrO7tGplDLUUf4I0W6sBXG4VzqipL6mt97
hIisobzWjY7JqhtwMCbb/4Fwu13NZHGY0CN0QoQfTSstErbclGtenN1HLEA8O2x6
ES5b5Mf5FZdkyNOEuYeXtI35qNl6u+UTJpul4jzHdh15M6Yl/m9bqeS2qOHzOWnG
fpQYuU49S5Elzw7stwuH3y1jJz3ndjkJiRyLiWDfgLH8Rf8b/SlgQHJcJKwotB7D
N5CFUMlT2A6qT/fwYXhz/3ytCCIBcOVs6VD1YcVws5iN/aeZkjsMoCNNU4qQLFsK
SralUw66OsU/NYLWbOe+HPysI+Mrq4Vs8CS4KeJxsok+14eh9/7s4VZvXfikf0mH
HkjmwV11QhRnDoS7KVQpci3vwjr726UANFppmFSlWTrweV5O4njYqx19O8rkmO5N
RyDL+ppYsKJBfyAWdBGca0AA7FjPLgSXSrCrAQ8NodMipPcqxplu6OttfAUr4kPI
VEI7Ru22NuDvpVeTEBDEElE1QzvXcbbWYIxm1dtXMAzcZ3Z3qtFSndVQy9Q1B/6w
Zf0J9Dl9jnKvfhSG8jZXN2qTKcjfQKh6mXd7dy93pAE5Ifjh7GqNew6CGYWo13uh
JHcxAzULg4SnAkSp4lO3p+DoRHHWo03VATatae+2qDjTzOTDOw21ZRJA5PVzL02E
Wr8ZnVlUPKE5YdrcfTVs2cWenpDI3KDi07GKTUBXjL0YEEzs1kJ89qXk5sLyLA/b
h8pUStQj/F5mg25k0zrNZXG0iNwEwae4xrovIxEwkFGY8RDn9diUq+bofeR+4sRq
gdVhT47CMrYy3A48SEZrPUQgGSR1/WFxQzAabeQDD120tmSbJDYUvxNCvzVZi0BQ
CmKmKJ+HAuMbDbNfSyunhdQ1GOsdAQXzJOpPvWQZE/oIW3iqUALOXFqXysG9rDpJ
ZGQLeOmXU6AETy8U/IS1OjAB0Cd4XVX7TkI48CIUerxiBN0BwEi9ViXWnDhs1EWC
54O0aggtmLELRQr2rxDVBcoIoMQXSYa/42EWksJJgG2K3end/PeLye0ymIU8rFNX
5nw7aCJuMyCfmX/bLcRNm3CpSEvjXkdr3cybF27YaY6SJ0ETf7PlZIskgtnS1h4d
FmJCPFwWJ3Y121MHS5/iX5BjSVDq102hDdGAZSu0uMSJK7rqB1hmQuFLZxBATzV7
RdjUt3nqy2XekxNM9iCQke+qZyVvSqgcVWn62JBbgpPzoJfsRxcBt708DoBm+i8+
8oVgSlxxOIRf/Ps7zHpIwpokHj3ZOaF8ZEzTPcFiqdOWK1rwdqaxwbGSkRtKAkNt
CQVqMEa8q5GpLfjzS3fbuXSEjEAzgtFmwTctGMdnJPlW7SANQ4VVpLHVoc5k5hlf
2ZLBoSpv7QU2sT2bcUx0kO9lvPAt+8RKipRhdQmEWYq57l0xRrMCX79qeXLnds6e
K2GBES89ksDO2oiLPLsO4ybbtmZ0iGt+pja3jJwOXhT5cLaD8JXtuuIWvak6GGGZ
aCh4eD8NnGomQ/+GdMByjFvEWu0dU0yLzsN/4+CFSTrr6PJEtFiRSCpp22sa6r/L
xwtzkPxM5uGE3iFfS7oN8yYaBe5Y3LGQp+figV8QHJhihog9AXnlL/msmsi+9rAH
iD5RfS+hdZAIfFH28ogN7olf/7clHvmuSR5Ot4R0ztz7fexTMWU6r0oaiyGvvFfB
Z/5LdpYObnCnEqn4yF1oZOMtHudqx4wntIIg670o1iafkET1OkI9Ina8WFSzUHNA
lyvkxhrj2dbyL2b+jmpFKI03Vbn7gHtv1p1BRGGZYWEMttrieHaVFW8Shl6kytTi
xJL9WUZgkIYY8Pzr5QVnr4trdqDGlYE3JySNETSyUHUsrVpXR+ZX5o/BQnfG2xb7
IwBJQs0uoYQdLQpCcY26OFWoORdvkFmWsLxmMoPPR/ROVFPT0SyoN2nNWPmbGfhJ
UBaGdOkT+mTaTmEfr8CCli9psO3E0MOhYGWFoWVqWvNLS1p6Lwoov1LNwa7h74Dc
bLeAymrZKiJ9rcpVGU3jjQFPglSEH+aVd6ymg4Ucf/uka/pTd8oHni+Lklqmu0Tc
OXnAZ5/DysH/+IqsQrFflU8il5mgHWy/nlAhKj6wIx5HVFcXW154wN0WboXpOxpO
vxjXlOq7ORq0HKzN3UpvhAn5Rq96x1+psgpThRR+ZH20S9CYe9yU3SJKRvyWTB5v
tR0/i4dtGtHK10fnaEZpBa20GzG6eJDN7SkSMtcm4cXq4xcsFevNCPwQrhsk35RL
ZK9TzVZBNGuMzkDxJj0T6Lm8XaNqQ4KCkJHYkQM3tyk96Gdrb0KhbuYnohIu0i2l
qWPN6TFkJiKS1NYbA2rDLILrWA5JxUTtg1IVCgr3fgvvkuEBNkaBawZVJSC6T/0p
4JF0D4HnucSj7acjzy40K+qWO7EnDK7W4kNrfy86k4nOqGf1FdZxnROuxv/LxVnY
ShPpnvUeLP8KxQwDVgmeI627Atr1krvRIyDy1eVVSCRjAB6Akyjzy1RL351LmzI6
ZMCcv7mU/L3V2zUsYIdja9ditUp6kY/KnhE9NBCL0GzHh24lyFYdE/xad4CQdw4D
tjxzi1Q+JGDCK+FBhCTgk4TLK6Ex/HDqVM4DdXScpyr8gCV9gHgnb79WIBQtQwT9
SIkbBJKNSOkZQnvlvnPwqjpEdYThZiuQJEL8mRix9SXOTHJrB/nOiA7GDB+KBDm2
8WBN5sUUYwBbYEIEyPgJRAbyype26sceZ8IX+zFzFfCK86r7Ci1pSmpwqDqhBmCP
HERT460IymrD1gLD/Fu37UW4yO9CcgY/QDteVGoPtJcpFyZzm5IF3PDDnbx1Xtcd
d7hv2+VVZ2+VA+5R8ZhF698kAviJ62F1kLlw1owubMZt+jsM1rH+sRuCSVKNs6s1
Z4TNqUh7Y5LxuF92cWlUOYlGqWAhR02o84AJt7iyrb6xThwWrnXyq45OygdVXdvd
+yKz21PTH+3TdwIo55s6Apf+rzOatFxp88TXihWoGnjbIkq5GFiqhyng3mzxeDFx
svkznCprtpqSi6cYceUR45g6FT8uxsz9OMWeklZah7tlyrygzfbXzlUgTyjRg3jF
uEo4jbUrUFoNIEgdb1hpfQyKu3OYMcodMKgAXNb8NztZyNesbAnI75ktlYcbOZzm
5Kte7g3ZrpZZwgpuJdKYd3GzQcpN98zXiZo926F6+x96xlutxeI+Nii1xjmpf2Zc
HXVcuyu/Md29unao44T4fLTWxLr7N0VR1TtYzmV3sg77iG7Vmat+DtqAb2OmSCf1
kE5XETnlJ2+QMqb/w1FO1zXQmZnGQBrf3GIs22LiKV2KDbDa5SFkHrOJ6VCkm3n4
FfjYXmf/b7TZE8OlRFvMVPp8nQ+6fslLzTC0k+jfJuq5JmGYAdqNQBnOH9LVPJT1
quODs3MUS4Pe1fgWTHWyHrojcT+jPaY8aBwxGmUlNG5oHjkwITXc5I+DL3d2OlG1
FRwVXn3QtF8t0f83sX0NOuah4hVPMDahvAevwZ1NRY+bE36wtScLvVqKwvkqsb2p
chP5RiNb19dmv5+xgvICQvwHb6PceRvArtIE3sWZaQu+xvC0FF4VjESfVKT9JbCb
LxVneU9pGTZP0J+CM7lvRRcG1k816G0Jl1q4Ig3f3Cog1PQs6z+tyDI0NMqkV15u
0K0V+bTJdMSHIJA+X+j9IRp1/0x/UGx+gHxGRgrNh00De0QjBuy2pqVgwEFRRt6t
Ua/YT+nlvzNOtX5JR5TtDthO/LzHvJCUKYa99N1ZBi0Sgd21338uR4w5VeX4oNYH
IUmeSkbCHA6jizjnQMWj5Zk4pyb+sTrJmdn8aVsbVJOz5WMOPKwlKLAZAxJQ57P6
js5hc0fzxFYym6JNTvz/EAZbs4zOCug1QDfc2bAt9iKuLUoi2+Ajb2FidVagnOSi
EvHqhBhF3m/qBvsbhNNvw8zEcXCjpIkt8QsTrbMi2P4kDVFGG2Syz4rhIFrFp9Ih
wIov3Dlv7tib3/bDeVBvb4/wTS4qniwpQaXlC3FRgaUaJN0JGmPYaJIAfHjj52kQ
48L71aROYnL7CDBxEbQgcftQUYhijJBq+RR1f+D4PKaI3Hn4wicFg/cl1Y+uQG0m
1rCegV4MUCurLzWyHd7mJQWg61YOQ908YUeIBC+ekvi+WNSXQFd0PbC9oxoHvf8P
/Ka51uY3wxStUYTJgT+ISWQ1reBtoZ21uPnCyBaxp0BBLHNa7Sxzn7t+6gbEkcNn
F3a+dLadGHLRamsG7yji3q7CZG4pQx1gvV8NUTAZBuUW7Kszxl1Pj7ezY5DGo13C
qY3qHWjlZ66IdOdha77fTEF2jLCrDYRWGNtcR12N4fU8ybBJTSnUD9y7m5H5rTQI
CAxrd9h9FmAEvJDQ7Bc6zrx8GTwmVwOsgk17nMjzHzvUZxmDbzAHTnmvwp8CeNW4
SYtnWMWLfv1VZ1J1iXYpbpCHgn9wH6yBY3wPoGFZP0A4GX4L4TwDsVTo7cYLbSgB
cfuP7HH8CZxgIcnpa5cvYvlGIS8+SzO/hLqHREA2awZF+SZLsEkNVAscpvf0iNAp
tw0mx4FojmRkeJ/atsvjNGDLzT5ofUBru0W05+Fwtm7QC7W6EsFeTrlkgeFEy19z
ExfB4lrsQM+euE2dlvR0X480XFO9TPOFahySAlzPXr40hC+wKrAOgDokttcS+LBr
c0prfNkpsZTNSBBFcliJ6V5UyVbY+JBjipSTVDvUg9N9zKsO0VaVRxnFuN5pGPXa
B7VMvMBDvpaki+KF7OYYayLden2QSynhRw5K16DME8OdGeFtWiZGODwJHmuLzCx9
7WZre+JUCc3YsiEkeKoghqGFrWg2kiOgJWDdHA1x9X1fAMBAq+7kUucVOIfUASnM
V3fy+jBbTTX0C2BJmOgz2iJ1SDrV94K3WIkQQlflWyx7/8jC8Ts8QTMbBzB2esh3
XbIv2VPdAnrVhWExnNQ9+/0UO+Pb+kfCsO/RpK1lgyGk1K5RE/emzTQmK/pV23QV
jrywvTI73xoDhIyNmIs6yIpEYC8bjqOe8S1HX6L1V3SxIn9N2nmJG2GU0TvabtX5
LPKQ1HqoJ2Izyj1XTWSSSnmjOVumtPvPKn+tG+JU+OnRT3xm2OUe/v7sC/iGrJmY
P869a8y1w3kY4mOXnFVThpprpB+F/VQjKolWqzMUK4h6hyNugVLtnf1VdsJol5yE
ZaZs8hvOEkUdpSmsAKk1DBsMnKHfSj/YtkrmWuKrcyt0GaHOo2xXvKsI1V2HHv45
e5secDn0ETE8N/NFvZZWoogwXQwPD/xfRuThH0uBB91Ef6n/jrdhtuvdfm6mTNjr
CMqTFwsyN3LuWGvzcvf/EwgVHDtILHidk6CRmy3DL1snFiobpfeYkzIXp/PmhtD0
92Oa+LHBBXWWiTtgNqB7NLZFshixcUHwkc3e1SAG+Xx3vLC72l8aNlCwag1woKhS
Lqva8jYs21UMWYPj9RtPHoVVWGhyII5GvXi+we7feOmJtXfvDOLkxMUtSfNUfBwS
WxbbF0UF+ezQqTSTECQCHx1RlRLny010sEnFyAdacLGOBbSG4ECbDgihXX/lxiL0
SzIrRrmnmKAGnWwawaUrVKESeaOAd4eMG2MXFziFy4L+Wig+kZegTaFHLAQaofBW
L/ynRhrzIbWEV8qsd2IJRGIgZBeMT5NubDSR7OGI2z2n+7b6RxoxREipIWFemEyM
H4PtbSSrVuJWNO5rCQ2Or/YWcOzPqgBLVi26GIyvGtXU9yhDroaGOTEvzjt225L/
y7PSbuXznQOFj6Kv6ZmojH9NRONFYkrFKfEinM6mb5okY1lppV5FqlgzIrpZpXO0
67Cbvyp4VEOnEJwHETyQ/cke9EZT1vtTFmCa5MqerEWOLpbGVCi7bcnSEmuYdoUv
ovf1gdv2+47jqmsWTW7QG6ZMIMIexQShCmYsY7IBh99mmDju4CVHkPkZr5hWuasm
GbWfv0lI+SzwbttIldClfmY4xF/QwGSV8nfiVrcLl5rEZYyTYTND3rjjPwSi1A4O
q6lCe0ZWfPdF9ELV9XmFSjuHLeP0Fh+VCEMyLP61cW6hsIhPWXFejapFoT+kUyyi
/K4BAkpBdHh+dMuDDFW1Qe9/VZ40kCaOwX8XxqUYSIxepkU70MJfY5aRHZxEuMUy
vJRvPFUp6UbKL5bQDyKoCjZyBoKRY1GBwgQzdIWVep1y2SeLXKMNHfKmUhHTS/jA
YX2hlSftHvZkiMMsGIDaZ+mdgBttCzIw8NxtP+x5p8HOz/SVj0racn9jw2BQ1oDo
vAgy/KJ/HMt6Wgnzbv2elXOi06r+qqyh39c5LB4J5m3mReXRnMRzQarKekdP2EEV
I6bIPUllVtgDDkhTm2d9bkHeSGH6QGryYPMR9dtTfWIEEKYjsIAjRXri4mdXFhxD
1t38TNHGYNy6VAFPU938nUs/Z7Vq+l62/OhPiPnSr5X2QHPqnZ/s0zQndhmdKcXa
QVywJrixrWO9MQXxT4IAx3MKj51s85An4OsA09qmKqGgzHyh2rV1HAuOtmmPs5Yw
l5qA51LhIGbUAUkfx60wAqEFe1fDVllhUcoCYKMIGwvpxjtZA7TbDvbClvTE1p1V
6p46RoL2gSt1RD7UfvnPGIcmIeAz9zJITY/JdY1fdW7MWv+z4/tdDDFKP3+/LpNf
49Hj6jtL8eQ0xLrMrZDS2vq0ojCFMUWK3pZS88Mc+elocyL0yY/N1ivSH6xt9qMu
67DP8Jeoex+g+qry8Fg7Powq8u17qHAPktMB5jX/j5mkuq3CXrdjLjHvHnUpyOMq
sjtBgHymTXvkTNPlvWmcdvf1TpFxjq4BMS8V2Ub1ss7uPjqEyMnOcMIZrZFecV1p
7zbGA6MHt2mIluL58o34x8mu3xgniTs0VRcrnoS8fcZ0q+tagIfdcJCSwNhS340t
Say75kXOm3JT0mWfs2zSJwHPqwrflAVQhBzRJOp3RurvRDh3IBHBAWEH6bsPZL+O
7kQ8cVlWv2TiJK89HqcZI60oI2iowmlkjKAQ3ndMS6YmuqiOnEcUJNFcWC17Dt7d
BimDxEQwg7XC87rk9EmiIw3RAU4sW3z+wBDYELAYoFIW839RVQEIUaBUGNhRkc3w
Am2g+gnnmotRr8eUB8VpKrgWXi0vMW5Mkb+DvrwSZgl4vUgLfVa2L5xCUc25RADf
da7fvqDG8Ko+nIKyeuGF1HtfzU6VNUngzTxUulTvuRM9K1uxYhz4QAdqwAh1XgXR
CEZ3NKk9RIz11ZUfvOEgeI4DePJ+iLYHuZKjq8sql18whxx0xTA3tVNJdOFVueYy
kF+vnsXwp+VAFP340qJ3j3KBRIC5SRNLsYVxzW1YxSky7RSofVWoXJzyguADqFSm
UySqBFheMdhpRWgxJhuGytLj9kDe/Kv0FAnif3OkPLDuByjj9TuDmfm8LruqjsFg
erA2H8EBRWcW6MSJf1D5ZuXLZDH/6gGq1LX/pdJitTMEOb4GEHUnrQ/cJw1YvlrG
Tms8md1hXt9ZP+YvYfz9Wm0nHW6NCYqPXRNax8J5ey5f2gB+4FKJso1pMEB2Kc3V
TJTPvyRMyalOdvrEmhxcNB8USym5iHdm0vus/6Pf2/+N82Tm8wAiWcBSWarFZo5X
LDEB4hAjDLtHFLNmJ8WEzKNbOTTfzgHqDOuyEsMa12SrcjWAmVVI14TJQ9YhT7KI
zCEUKhowPtDiGelp9fC6ezKfftNWxiql88+jpsiUIY/Wfc6YF1clmD5rj3ywAi4s
+5/5sIgn2sUmiz9eIiBYUYfO/Y4szmiWoVmSL2PYSpqYA1xCbYxo1vI5kzd/bAl5
+pLFpcPs5zCrjDbffS6shppWICD5fvNxCtxV7ISwWiJn9xZHBI2EhEwyz3R77c3s
W6j6oY50rhJKdbYh7QLON8MNSG7g6UqWNKYPYZouKgch3ohAyDOjwdN6VTzfyWeX
IDhrab9YKD3j5isp9wEEbliHyAeKx4wpKOGq78LlxUB/MYV36Cboilw60AxW0vYr
nuIdKKw2eh2TstWW2EscA4RYTd8GnFvtd78eMF7Xx+SagxVV0Phyf0Y7XvkHGmYE
b0rJUVrUqaqoZvAKDyi/uHIUYxNxZLz6XEHGtkQNQ2fgbIdyavjLspq7vjKv0jC5
ekG/Vi2Hy9Mob7WKTvxy4Ja+/EQcj0dpWJ4duVlWLn4TZGE/GTe8MFhvNjRak6NC
VemWlysxF4MybUj+ZdMSIFrXUiZ7oinGqRPF5kJgnrCEpPzzI61mFH5N+lz7XYH3
INU+V2MdHDCgPdYbNFqf6m5nCZ8VrqH2IQOF1Z5cbxKmdQOyhFf9Q6jTs13sGgdk
Nt10QnENauKuUinE3lk0imbqBUOdLfWMn8x6zr6A4x0qNrWBM4c+6RFKTQEvCVRd
Rg2/iKItLWIbe90YJKNBNhX+U0Pm0wnyevOydgvzJ7PIeZt+HVTo90Ugyy4n7ypm
kH1b0OKOOHbdfHiZojhfVuGxPtoYC6Np6la3RIB1AaVDplP1L/gSaXVz1m1COV76
NCtQPCe38TRBpGKPwtAYB9gYvDQxyJGpcPLWgHrUh3cM0qfVyNMI3GJWutTekMBM
Fuk2x7fTuEnfP9h0L67Y9UDzXvPt9Exj2n6SKcRXCD/jlp9/3aKkgQTv/FIFpX7C
WwQXk6a57pN3HIP3M4FChIEL2sFLKBFeFtlBo4upaM/v45GXpFcXSWDoRAEUqSxZ
ehI1MRh1ox+F4q3cpg6tt4VY6aokUvufnh+3DV30CC73tibG2PNQAZhKEJaS+PD+
L7uD1H46cYbSORe/KVDu0EvEZgkNZu3DSojJYbLgv9nBTN7jGZitEoAxiVrUsHLt
SUg2VpH28+BmIm574Jzus6fOgImG2DuDBc+Moat71wRfuDxnnMPXU0TGssPYLikT
uxWf2wkK1OxNoIwo9w/hxMh9prC4QINDhErZEZnR0n9f9tyK5P37OqD1kmOJxHRl
GsDN2lJwBh+sJlL/9b8KNNcLw9hgIXovET0eIDQu49z5+DEf3H2JPbACSbmvBxmz
04dxQSqQTKF02X52Xn9pxNxR1CDG5VtALzIzMATXnp5WxzFhF8Al3JFPWiZ25uoz
7lllM6ifJrEqbBwyeCE5L96Got7CFtnMhEuwF9xlZLVnVcIdERnxO7Q6ehETzRdE
pXuNXB79p8yovFvtsqKiN873ogF4FdH8/FGw9VMV5vxiet+G5SjpKVyQZNLLLFOo
GbjAbfF40vYBWwsXca+SJ7MNn2laeJBVElDqXvoVdTSbHNubdIg7GoS7FL/WgKYE
LImFV6JJ8MiSexY2NyW50tyCEJO/xQjYq68ZlbdofiWKBaRyyLyH0jWuJz6hOIhF
V1o+tGgQ7oSjBTFO8yDfBC8sl4RKH5pwYOdFzbir2GEIoYQbc4zEWqcLtP7gvqid
6Uk4eLwOEqF6HOWacgOPUcEYl+aEtlHaXgX/K/RLFgCEmGLdp0FlX5n5nkaRqbO7
dEuF4MbVxcytS9jOEAKTDtd4jx0ARKXw6C37PyB7I/1nSbppgVHPNRXbHNzmKn9m
XLdYNg3NozT5TZj3jMAnWIBqrHSQpcKlyamjSngITpPDdYOCfa8mOR2WzSouTMVn
udkX7mj+AnB0R1+xWbzDvbhmKEIgX42qT+8iDRhCuaYfV2OPALhoS72bGxj8whQN
6tsqlKlMgdapc7nX7dP3F1K4Q3/1Fu8DD38AWHNagT+bm+pO3O0sAgjZ0KzpDp78
zxoVj5uBLGDkBddGtcUSrI2o31mXf/5Wiitd8adk+BFAU4Ob4vUNLdnobqfTHFz4
gHyGsB/lWPnX8wsfPA3IxC37T0Wip5HdGN0PDc9pgWaxbnm0nyBQWSwdHhx7f5FZ
Lobl24FTBBaVizwQwL3fusFECMM3NKzmncBQGsYBzKgChKbC8jL+lAk8jhdUpfSV
Of/LmJNAJtehCxciZkeFNtKjBj9V0kBSHc8/1GL/irUserZlXndNmyIqlE9AJO53
M+zX2gs0xNvhiDC4Qme+KX/7p5JVO05x5K7XtLB4/259wjkN8gbe8TTNKCNU9UYw
8YKtBIa8fT5+ipiMEYdtKpDHgc53kpyXNGnSvRruqGuPeAHaiD29umXfG9W9UdDW
hpn6bvvpkCLFSgMUymZYYUJjqI2FkecznMrbP++41wDJ0wV4923vFEdnBxfS+Q04
f0JCIAZAU52QXzmwTNliw3s4P6H2SmW2VOUuPn30umKGY6PaHDxFYHCjSX2lgYe/
kGZpdxKCBytKiECXzx0dq5g1qFr+q5e1+5EX+4ssONfjsJd31p9ZRY2LnPh2mHI2
PO/A45bMdIWxad9KHxnMldHqP8qu69sucA8EPImLB8ukoHr7YG7H3dj2wPiA1UHO
NK/gc4ovR/2jWrZBUVtct43GG2f3kveN8TN7ouyZYGZ65KWFZq0aK0F9XAjaOqda
5wC4VCpDXjVfuzh2aG6Rjlcu+gSE4qdJMVPQdTRhzHsw9xvnr3+nQPjOhs9eARCC
fZCzZegK5yBA+jFHGC1wPP1uKTZy6G6vfTsZ0iZkwzJXT2hvg5Nqpc0HmyS/BKU6
LTlmKEsx3KITCFw5LNL6Vt+VTzHv/OHv9VIe2M4i0r6Gh7xYQ96Q9/seMHhZqziF
ehyXzrJPw99UiqkLBDSvpQTYCOnIE51T4aVVJQm3FQ+5i5fPEH1dcE1e6mf7jkKl
liY5zW3HEV3d0orFX0eiQ/jOouNYTomqCJt79Ochv4MLo4FMd36fBZvodBt+58wU
QV8RO43+eNsMjfDrQA41aaWm2iYRdxNdfhdT2bnO5gySaVqdx4QUjPEUAc1M1avQ
Bpl4B/MI5lpEkaS/Y1Cc6NdQjscdzDZLLZuR+SzwlGlYwZf4Tmzyqgc13sCRhHw/
oZNjr7Qf4sSBthKHlg2TKcJSqOdWdDDjtJtBS80eQAdriXnP7r0b4WLMAZljIqTx
w04DjGB9eo3IRcczt/o6b9CRU4IhzYsVGxNORKJMMAnFLkrXlFmdH9338QseYRKt
8Pp9LCY9AmAPhPZ22xk76QYR2ZKTIEVIp5AwSFHjWT129B9ZtQjnvz9xcbBB56su
F5HhANWz7qf6Ff93olOeQa8+qtwcd1z4Q1Jjoko8ZZtuQaDRCB0npHBNN8v42fQz
JAcvOQ/00O+U4GxbFUpHvuVGqrUAWLu+xnaqwn4LcuFwk1nmOAaAif9UnYwQ2FhI
mGymFi8Hyj7cC9qGeE9wQnzb3p734evbafepfkDcMpZZ80ts9A2xWQyirh7TahLN
1yxovq8dV/VRB1Yp/9Jc77DhyyGF+ZkUespIGy8WrOENtfFskab3IqjtaGkhI0Jg
aFC4kK6CuWZ8gVfgt5kThoY9qC/fQyaxTMcoEydE/Jy7HZMxoGKuK5TNP+slioy2
vjSKKc2EGoFcHIlBy202UC+mdELV3ZuZQz4s0bhtTqAyW7Bhf2QH1j17A13OJ9ID
SU6dj1VjZWKek6wlcV805YpCeNGQ1HYWaRhGNOqHK4aOreJdD3jG+Ds31KR+Odjg
WJ4GBxFwGA1Yxy0bhGkO9yVoJNWuBJgbDUtbPIzCZB7gr3Q6mgFMeJcjxI2FyUTr
AURaolJeAzbFXlg3nJEsxX5PHgxY9vZFQCQ+WHPOIxlkmBZBqFBbv6LY9Emwx2Gl
0zN1Rcm7umq2y0SBpZcSPNXpkpRFWXIELRPi4HNO40NZtx3dbasTlJ2XlFpRkrow
BU6JoW+/QA8s0TSnhb+G6gT57G5oNMcaHUEPKTfdCKsKL0+2Mlgk/hI/qIUnVQoj
fDat9+88ngWfksg+y0ke6da9Hk3yErZg2z0i7JPidhZvVffKP+KFDiLxDydL4dWe
+uFqVQ7tkcschjmVvjjAAvCrD1v3RtaMU546NRZ0eajB5RnDByQ7cY8TfAMHjGyB
qtb/acAmJwXQdUBZusMSgnNlRGOuEYAoTfOE7NPZPfxl5m5TW4mkbAqJ8aoaPA+z
TUzmU47Ihhm94yjDoJHcR8/G02uE9YmGiDA3pBBtrIHMAIie2+iRGdWZfpuPar0w
njhblqC4qO4SKDhdgE8oM0CNtcIGLxYrMooJzYfTrumVyIgwlLvLQ4yyUA+u6B5v
x3mFn5hAC9IRl05cRA88pfkKIJ0GHgVEdBo+h79VGWZ71F01oS/zzIST47BXFOkb
HWGO/7cOdiuL1EWORCTDRyb4z56grFQd9YKtmQdyyN+Zww07T6HjsHT6eP6nZ2v2
+G2kUKOxeFJ7xjtpSdIhLa4Dl/mczqYA+/6YJc+qESmkTo6FZXUFLNRAa9RiGO2m
JGljhFDuRMoKSs7En8lrEstASQ3gU/XCP27K7zFAflN0SzEXsi+ms1nXBuF2stgh
MNbztTBNp6kKb1I4TFbwpMIbZKtf7eT6gTzKlDwTI+6EiHzBNWcysr6pQq7cvnZ2
aG5d0at4SjYwk70Gc7BIfdS1QgBjBtUvSfeWbifI6i1ayepziKh6dCiyewQqKRlA
7EVGybZLAjZt3DZJPlZHF37ezUZiaoAeLajr9UAGazpl7lHNLcrokPfg5eZOywj0
BdVHe1AAEydzCE41zWzMunkTj/hqVfigrF2E9FONUgJ4KwnumZvsBMFQKEbcP8Sr
8STmRvnObngc58MfKgAfkuYVUFZc0QA51Ymqj1Ffzng6ze7Fm91GOS2GUu8qbS6d
ydJ+9xgoq87bIYoSWW3J4MF9bs0pAjR0BHmtarVxgemeIQ39nzPTikBvKHyk9m7z
XRtQiSpUIRMr2nFgnz3sgza4jo9/xT6sv2jKUKcB+SELOW+LBH90wf+LO2ApINgx
HTf6IHAjQUwpIhYolzX2+EPbP7BfHZm1DLCJahxrWc3j/VLB0ccTfFS0ecwQIKKY
WIveP9247MxuDuZWDhQF187tKanMH6jBhr/RKMcSpBXpM+blPWcFfK5eOGunktYe
2WPg8gZC88hSC07w01RH6+rVFkYC73MueyHKq8nbn9xkjOe6exGfBezP74FPQ46N
3uQCriEvpHPzLS0WRqow3qoB90EeHZx129zFH9KX3wZv8v4HgnyR6EouD08og0Lm
tJmAjO3MXLYt7G8Xy3UUPc33bRbUana+1YZNKwEP1jG5z1QN+JQC7jtIotz+RiPa
zl1wG5D7DqqpSgzbzdEWY3Y5L58PADOSaKW2kXvKbhgJrGmLqi2WDgtgWgy9oWUJ
bkP3ZkeSI6I5tv2+GckC9M9j2qkzz7nU/3GEtFuNi/QBB6HyIbHSLt6QX5MBxDxO
EPlv3ulemMWZ7R3f2y3MkfcJAwp2cS1bOCWpwfNcr2eIvGW/8krXpr1VkHt7hz0Y
PtHlucQuYsjLZrpdJU+J3ozdIjpoIcBg/dL33dEdEG54YcqN/JNtZYPaE5e967Xk
lgu2laaM3i91Fa+7bOJQioFu9U4l047LJYyy6UAfT0xPG7SWESI+phhJKL6Sk8Vc
O7v9vYkmHDBH1/jDpg+tM9DxZoyiZNoE704ASu6KQtoBv5t/3OF6PBV/82WJIwlU
RwX3eNZj5/78KZGo/B2tUY9dG2WgUrhYlvrM5+Gn3+PSfwEnz4uL0o0dN+OIc9Kn
Zd2y233ZXrvs/Qt3z9RQRRV3npUWAepN3TU8RYp1BJyfHAQOXGyq13ssI2FFrN7V
Gsyxu9/ui0JRf3xU4reLOgtGO/3BJpuioJYh9dlB7x/ok+l2ydw83J9GIx5sRP9Y
okOOVo7cetwWyBV7VTZ0FCEqFOMJdn21xex2L/py8+0I28cVmjEexMG00BpW2jfV
jTVD3iGhc9rmMAHdDIT/AGQtQ/xsAbbV1vVRgE8VWY8CBzqQcoHOD0IbIXDGpLUv
rX7Pr22gBS2TZW9KxeBioResGixJdT2BOuJR4cRAvlfDzsTLdhS2WuilZheaJqRi
w+j6SIe6pkj9wngnVK4ZDIh5+2jgriNZhKp50s5d8+EY1aGwhmgb4gUfYZdGFfjV
r/9I725ByE30GkIxTdJBAFLZAQ1+t9bGqYgNhem2ltgc54xeB3JHs47IcWbpm6jo
j4GyoRz1dfybZVvYefsqDUUqe3P60QpyY8GP///4nUQ98yLb8EUzIcMVe574QAZH
VNCbHAZOpShpln0Gnh1Wu0xhiapFWVc4wg25ydpyMVgmCB403uz2i1BbXjKvi9ay
FSBvfX3lILBrDfLS0RzLlUgwqxIadNn52nDxUWGoEreEykAuejPabcV7iKhOcOK0
23nwgjSI19jjgJuFAjwlG6iJBAAxb60vJ5YYqGOFT9TYzKC1ZE93IPVJE0BDj3cz
/d/5Y7dAGOzqvremwg+BUba+kpjOjxIhYw0xS2Hc+KV65Laq8+pMoolCPieF87Fs
KnQH89rSVPvpA7Bw3NeTJrEWEDgbvw1sV7d/KYPDk9Yw/k6Kq55fFuSYeNagU1AN
K/EOFguIGL/yVFn8cZ2DoEb3jZk5Gcj86AEcltQZW3SX8lmp8DiSnQoeWsU7p6Dl
QONB2njxZPr02mI+xG+bmxLCrjWSK2c4ZhhbA1zH5HmMHBk7rtli8CNnjjYq3ZH9
4D/fC+Z9YMVOiMlSSfGsx9rY4X1GuSmK042k1UzEnw0fP8hlwdAvXPRVbzLpgW5z
movK6unhi+uiDydxthtV1dtG0liTCDb7P0MY+FiRQP5dbvgyuzN3EEmK0fuf2Sdy
AkGT12uiLNCtJzd3qRQdHsrNZacyEDXxLXDpYw2HhOXP3+c4n3D5Ges1SMYtGiQO
V5DG1a4jKHNiOA/ydqXAtUSGpz93PnLtGUw/fbGjs0cRXDOsSM/YolzRqCSNbm8w
95s9wH7OjtunzO2TbmT+oj91fZo/pFWQpMCAmChtlFOupkgJrCPy9FZRv3rYN0UV
JU8vHP9OW2zjDrE/plcilo3qv9MXVscoaImVVf2M3zsyufz97By7d+rR9vLDvUvG
Lklp/Z8UQTt6cMCNwAAbWCuENFTYCflyPuIrqVMCOYK0J4KCwJg76woulnvtLgQ5
W8xM0m/AXBdh5KtgQrYWO2uUf6Av61ZYNpGwYUicHzT9fXsIinWvQOmPHB86CF04
hksJ/GClxonVHFQHQmoY7H0pUFDyXDgYp1J8DHDGXPEEdAu5GLsZKmCqLyFE6CN1
vGnOnn9T3ishhAxuNoxD79Zb7xoro0/oEuI0K9CVS2Y7Apef++bKN26l0Je/otQb
XXecVL0IxNXwFd9iHtK7FtNDuwTLDVtrWq0cfoMQJmM+qqdvYuXS4m/es0CZnL4R
vBI4jhuVL28b5Eo6lvGyEDsAjn/F/gxDcMFD0VYopNTbzg5fGX2h5yEoeEwv42+J
lCbb8/GWf3ChM9jjq8j7tsg1bPcVkHQX3RvkYBrHs36pk/HeAwuaNBnD/CQE9xRD
IUx+jtm1dEIrdBJHH9PXcLcVVfFSsuU5coPyd9z0g8It8S2fFnBbYO6At7DJ0ZaC
1fgWzBptLNdQuNtCdAc4IrGLWocinW1xjK570Gkprz0F/L3ZI9DHFPfIgaU2VARC
5uGpPp9ho+hXuznl3DVxd0xqIul8jVvEzxcGfOZyZfGKXMvxu5O2Vjf9nWViMGvV
qqzc1jF3lYrDneEm8Cr+EVjOZv0ZP4rVsGZMtTLCgFszoJUUKADnupL6xa6BEdDV
BS3uJ06DOGsxjy238KISC/WWs0YKAMch2iKqZ9CXjx6MeeBiRoogBx0H1QuZlq7O
k8c2UX1bAyvvQdMAWuhYM+vBXkLVExfwR9IdGwuTkSFgBamxTB9A3mM4Xz2DeDjr
Nw5B8wJjT9Z29zmMTjMKJTmZOotUujDobaG8RgNCocMxATtqH+mcxiN2S0cwvh6I
mqDXaCxplDV3qnwuwbDIN1lKa+2EjgdMNoXEJQphCV0XrKb1von2kDZgZS+7bp20
8TaOv49n8/KuaY4y2eC3g5uuhAlLYl7ExU5elYkj6ykMdjiVW8vlePtNCnmwQDcf
c7icn7POpKCSFuJ2MRavBOG1esaVodYXfRKv1XnSAehzNaoZefFRZsM6Xyfkqxa9
rEqpy81IsbXxdUE6yHQkdsNmePJS3K8M5hMm3runr/bfSVzQNnOOk4XwGV6cZZma
CIqCSazziV93Zx5PF0gPqS3uvYVFQQMqCYs+uI4nOfL4cdCo1x9Zsp//82gD2xsR
F0ZaYHkOLLGpcZ3rTJKPHoIdoLhDDSjBLwt1AvzeHRbvuiKKSzA9B9bmw62T560M
jZpcc59V4hSnoJ3Si8DFQGsi39+8bjaop9swPLnf6TBJgQiM5SQ3kMU1jxXoNVzh
EsF6u7n50DadmzNy2jR0YrH855Cuwepc+UaHyrYKUK5OIkPfyskChZRgnZfO5sp5
rDL/86xtxwJYYTdLU8HUwxWslmnIBBc7kVtqeWPrx9nfREtcOC2+xsfjyMZ0XyLR
YQNfKPlFMgDK2iYyiulqFWve9mdaP7zdXiRlC8x5+VnFa+D2Ewwp2ZlPvm3iqjHT
PKOYDhAZNxYR/lO8hKQ4MqkA68l7S6SpgV8hBjoO1lNwAOx+AxkFr+PumSiHDEXQ
QgifnjOgcN15OqK+R9/vZlxzmGEYhw2xTk4Y96ME365sRoy9GdJ2hu3L794SXWfM
AqBUlw6MYEP1HmNvwv838C960ZTWDCtxaGAbxkXAOoZZiD85xuk+zaRGUbpETVCX
KFWcRUp+HZeh8DiPTbQvS8aCM5mDWVZIMUHuSYlotT3AK2tM8lLPvmW9HxcetzQJ
79t7V6QoxpUr+3d0kK80Ao5FfOmxJBamlDUnrhnVPQTdp7a2yjE6kcvYahrnPRLM
UeAO2cNbZaCEcgT9lcflhsVxmvdcKOzNqIeK+CPh6iK8w1J+TR+GLRts/tj0bfqH
cWI07mpZcHh8VQlwKudPGARrpWLW4uIJQXdwaoPS1n8kycLhqnCvO1Mru7lfXcFb
U9hXqVLyGjl3OI61nPe2e+7vRgdlQ/mT3XRXGRnRwtphjkzSBcpv8HHYv1+yr80I
jlkfiQ7W9pXP7LgnxW5CSWg5K/q8gs//bcR8CFGUPk2QuzRO8j9LRmvUoxWQtaba
m3PFvgiC6ESLfWTV+DXf3+Q19VZAk86/KFJHq/3oVB/Eq8yUntTj0KKdceqvG317
vzvKk+HEWp1Jxg3lNcpv5mRIH0nBn1ffMR1F+Q/kW6YZ07AexZwoGGYt6c1ZMeRd
ojALGdUvnulEtpORH8dXWYzb/YzrACiH6zLqVKWfteEvovvyId+czaf9ov9DrXPe
5aqm9NzRhn+SnokDSwR0ZwG3YaOO08F49bQiGb69EY8+MYAuMyCSmNp42ZTbCsHh
0Kt/YeVdYIXfv2RRVN41U1vaxkLEs3WfVrCNfFK1rA4FwCn/wr/ojZLIr9XrriEr
MnVfrCJl/BiMnnzddSTIlfQ2WFbW9+Djhb73dSxa9DUze0ADysTWLtXXrZSrWVLD
37ML+ASvs3epACNwl3KxoKyc6lIGwTNg8taVW4JqKxq0AsA1UeDC5Sr9JAul+8nN
hRIjOakCuikB/pEfSlIFat18EOHniTu84+lNrYz4S/P3OfGD3/5f28UWWNpEzrBU
HnX/jKbJvyHwXRckNo9f0njnrapx9NOjRO9AeGxsFJKyUoS90nYDTf6M+7zjxohO
kepJJQkzvk7Qz33i2fguzXYGxGJ1sUFVev2oy1sUkrqsk9fiydyd8ocKv/q3IMRg
wuOWYCepxWNs61Gvm8XP5/B6rRrwHbWc8sJqxGK9d91rbM6BH91qupqgD6wqkz3N
rnf95R+cJ6HK78J04QOHK7C7OqyTGN0OUFxZ9sWrT84P8OKmcyUGX8CQ5Rlz9Q3G
L8skOJ4BETN/BSEv4tmIIpi2PwRXbHq7CsbUbVljSZKCbAtKKa1n53xgAEfwOHuZ
MzgDBg3lCn3p515zN117nC+n0nWUHDfl+yyEpdxwJhZ7P9zTPvEOfW/j+JQeIIXP
cs7EMZdtdj/FKmnGB3mBmrOYVb45QG5NlEwstIa8vJdrhTwg31E6G4f5cIJ7sbxm
jBKK1bJNuM3ahjzGF5RWoH3GaaYc1/aUXUmgISy3ivsA8Mk39q8tMUwpFhAjLb9E
qwU2WIgsyoSQsS0imnDfDA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
A1ObKt98iLHVEgnuaFZ1eQLAFWrEwzdblrhJa6pUiKFyau6GvjMzTdhsaSBiLk4Y
492tGLftMiIyAF0+R3he8fANIKu2RjaO0IplRKEICwnghZFKVj563lVzcD9O9IQZ
X8UzkF2H9f1bmbUGkVHytIe9ZA2P2AnrAssOLBQuLTSrSYh4UH4MMttXLo4Gr6wl
b+js02B5OuWjORqNNfBpbyS3ukZDAem/Xaha80cbyurG9pbqKvFCM/1rBqOieGUp
/ChFdAkDWigqayzXi+BhQFcEGZPjit80cOkcEtCtqnQ0NAhyvgAr1TjXFeskuqSO
jVVL099dsY6w2m2BP8w3eg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 19328 )
`pragma protect data_block
tJJ8UE2TECruXT5oOOApU4cmi6lvdEyUfWEywFOyrC9GsMAMvpSzE7u2lRoiO31V
aYQQOFNdd1CKdOE2S+ksqNHmgn59Pl4gT9FIPeSOLU6wwd2VXYUC9sLCRumb6qL0
xraPdnm8GrKuhqw+N5/FnUccAUdjThgE141LK+sVHAAuDEBDJiGWxGGUTJoxADEu
+K1Z7Sot36nv9Oi1T2cYxmTq6ZxnfzRZUs30Qdq4Ddsbbg2NGe6OvEyk4z+BYjRw
su9gtKhwVeImVSSC6zZaB+Cwsys8P+o6WzQNLK9kqeeh9GH+9S+KQtIdQAfu9A+5
LMULc/F9m54YbGttbTzZ3VzXer5YRO7xqkopJavxyXUqA4+rvt9uDrdcCpj8Xrer
ZK0ESAA9kwZ16xArl6DPFjAQqYaZM/whMtEivXqCyclsDQn8WPSQ/uCNEEj0vTE/
m81d24PqU+yr7A0S8vzh3fvEidVoStEuUO8HoyvcqCzKhpDt/rV/jY/Gkyu+XUc5
HxZ7QSs84bgdapJ7x/2fucA0m5TBzhpCIL/Kfr5yVnaA6/L61yMKvq1kpBSvl9ET
a9wf/Q365vQ0qcVXjoftDaHXKtwNDaP0lu84kLYWvPjP2LPmeDhcpOB6Is7gJ+Vf
Du/IC0kIYXJMWre8qAPD9iuHD9A8GDa9bBkgIZmGd9MHdB58gS2QOuy0cWWWGdoL
KDsEv/UFjpdPTgZWar/5ad6x5ecMhodr7yZ75JhWuiX9WrBMyu1hR6g5TimDVnBa
O8Fu3dYB80TboGN3B9TEIi+KpFGiMp+re4SE1//aBa1ldCvQQizeceQ+bmerG6X7
Fbl9DyXmfRBq1/o9uQP/tzHCBUnVrKxUqcrceK8KEa6rrGGtzPtydbqpiBp39VmU
JtbJuyjOXV714y7G6xvHwDVt+nMz30eJSixVAXBK0bRk5U6IoINDf9+5RTsqVT/Y
6DEsm8gmcK7gCSvn+atgJ/SBhmBDdwVZuPV8EwruA259u5zfOU1LpXoahf7XFH3E
g2VKm1B8mgf1ejGF6BwNvkTDXr+h8iluox+jrFd/iBOMK7nITT1xA2WYM1xnwuoR
JZgNYrBHI46AwZaKyG2utAnVLTGdZ1PhuspsA9zxcqOPaeEeGKJL38EwWARJmg5m
MzUblCg7mGvbp/8KInwSEeQJDbtvIJPWUlzwKqgvP/mmlmxeM3mJpDB+ihpivUQv
GtwjPu0NI1h+geVG1eGcncSxFytg+BjefIkDt5SotcipX96ir2Fh7ZzZs686ii3O
tgBkBRJNISz3lYUX8vLNOuw5gERnyFgP+ls7dCe+Sv9ccthlrJiaCt6CBEw8oDW2
+5G0V12sFNs0INkCkZYIINYsXPr8phfEF05FiA9bsW1a295F/Oz0hYNQ/2qBQrpo
qSZ24iipu0GgTZ9+nGnstwoxPpJwrin0bMuVfrZ2MY9IQqLhm1R+DQP0jHxVyNkr
tSuT8rHwyzkE14SddwJ/clgUN1Ra6qRzcyiMXWXtow5xsoQR+t6KilmRrukfcRJb
UtPb4tlGKKoMg2cl65IVzJxw8oZp/NiIHPiOn48CFGk//B/pnzor1egLQAIgqU3p
omDu+tn+/skExuSuJW9kBf05hKT9nmfpdipGVFKzxMoSY/0BFyKwOdHOmwrKNsFw
35wABsn5vqWa9DL7Slg+T//bYbQ2I4VwWKT/vbUKYGfzx/e8bMFt7wqSuz5xonos
oyeeqJyLyLJoFRF5gzZq/hfiekGQyoGh3mnYR6CTB2r1Jf4YczQZCRiyP4n4eWuT
UTn0c3xf+Y76q/thqDgpHfPsi4E8ImRhBLvzncW+pX7ywhxyRl+dEVulwmro0YaY
TerGWzNirSVz2LEiiGIPbnM0OEM805ye3g12K7O9AC6kLdShMOgCu9NrQV7zEjRu
QHvEnSjGZDAUkk1uwt+vJyTRvnG3JUqot1IZ2eaG+mQsb1vkuBu9NvUBJV3wPJ4y
UBn+ydU9ykNf7sk4S7sxt+11hxovm7pQ/j2BgtuVS7k4ZCpYKa5Q6V0VyoZNCeUv
2B0AVZg6s7DFONhM3XRN50gqjHpaSzEpcByPELlEzmWw1oi8bhKs1fsGSU1BoI1P
VmIABJRPoTssjriNor7x65NmQbBC03iprd0lZuSWDRjubyJto58tQGySS/WKbdVH
439w87WUBolj6GozIj1+D4UcskWcIXToGp/zTq0dKVKxfuISjE1T+/S9WLPKjjyg
e8YXfR289dh+pVNndLV+xo2WFcq6SPj/3AzE6MNwuEmpQiq3WN6e2H7Zf5rYBvRQ
0bWgIbN2DNK4UOETPA2GsQILdLcnxqPT8JJ6mhBaiq7w0fsk3/j+cDShgyS0lHp7
UcDDAwxHuJ+3ImKtSNCV9xfwYSsiTiGJrezi9+0ED3Q1EeCkxW2rqb+klTp8KGOW
IV5kRySqZWgeb91yqEpEYfgUoMDoCBYvoai+H+46LvDey60Mk+IApzMWWmvYKdqY
mlBBu2OeBuL5rixO12WeIiUfUdD6QAT6K807Ahn/BBJRbWL2Q+ex6coJ2AKQqvhp
7gVcpM3230hdAFrAurQnf+z/GBXs0Xo3BTMV7Qcpz5degCs2Df5hj9OTcnyoPJDc
cHETlechr+blFqNbgaHvXVhYGWWDaIK2QSUB5YYDUCtsQSREzKYwjOwhys9LQYZD
TrqL9d7h3ReKDcpNtRkqqVe233LLVhKVUwgS3UPSd9soQLA9sT3EiopsEdDP6UJF
o5Y2YliYp0o0wrLCF9y59xhBj9oZGw8DXY4TCN6n0yGG7ul4QOnwKK4d711tzayq
+fePSFBLHF/9dlg3i5vN21co3+efkANbx9Z3EJglD+RELl/kHMZFE0nF3hfp37G+
MDBSLAAoazd6b1RUw8WT9ejolylqDMm0nyvcQD7RbQxrvUJ/SppCEGZWyG7YO+lK
eJmLL7+zrVHcWFXAvaUIT/YJyoKeeF5UWtcaHrkhaoAnqeXz8PmaOrFd/8g+9j73
UAGs1QAAj/wuAXSL5N91fwSLrUOgnA5de39rySbc96WwEeFCz71zsRU0A3URtDhf
Xn0lboBayYVCQTjqh2FGu6Ig3RLyoOEJ0niL3jc5mEPTW38ObCAcTM4cv8HHBwEX
UwwTVrSx3ntr5zki0aL/RyVV56bE+WlTY9R9gkSc+u8UO5hZXBe+XRbY1x6LfTUT
2xDW3xn5xdVfokXiAZeGis8OCUWbYu5aO/hCc4gZBR1jPCEZKs9x1wjl5EIr3EV8
p/VtuUacSUtmNvwDV5EmmX9khxlH5hqTGLcy/nfAkaJ8O95uO5/e4Vla8CPmUMgh
ZYwjHASPAUPqqjd6rvuCy0+9ETT8lfopI1K7CAyFFldIPBs07zGXMjlsfJYKHKy4
9KE1OF4D16LIV+/fMGEuFAvOIS20e0ViMeqx0spH3xlZCfaXil3Ukhyp7H+VAuJv
LH4Ykq48J+LnvxWpGCMxdSxlgsR1xM89yBg0P+yj2llVxGw5wK7M+rOEG+VDDRyG
DveQYeajhM9MVQMcyy8QLQ0zSducRYCaEhA5gOsFmGEDS1I1SR4c2J8njBn+ssV0
Zs0a/jWKDnhHVbav4qZFyytiie1mTpyjCje4tRbm9R71dpJ/jaOUhGhXb3yIrscq
5o6PDSz9AivxYx1+W2d2wwDJLJAp+xqnZqMw/ZOSQ07jOEJWa4rGYpc+TIySmSj+
1UolXrjFEPYJFPjvrGbE9Hb/KbTVuKUxR7lXNXQzK+/FOYeK8Q6tNoZSJeV43NoK
u9tCX0sxVMPcTkfVw9h09yj/HeM/G0EvrSHzCnebTr5gvjIeDPopgISxVaHmHLR4
h1Dodz0Ecyrpl2SQYa4zF0xd/Uplwov3Z1j5E5PaJ6Eeo7gLRXkryUJvAF/wdCCt
tOX9jGepzsQmGXR7Dyo0SqtvIiGsc65b58/AAxXcroN7fFEmmr35LTlk7zQkwrqF
rENcT/Im9sESocSqdJyKdHH/JTrfhFgTi5Uq71QC/NN7+wIHCzXcVxoZCiQ1ufgz
fmXAwJE2X7eKAzfyf7cwQaqv92TQIyzSMICUw/AInNa+WehVdsjnp8E3QCbC9xG+
75mbMHOlEOhgQO6P+wQ6pJAhxEI3igbSS7cnbnnVpr9x44CP9+13tMLQ6YXy4Laa
rzvideAhCFELsCVZthn6d7kCXPZ2xOEGYckqTGSVzfFH6gHn1hzAYWIUd9G5gPu/
fivA04pB4V1wfKpwPRY7IaFyTymjDVbIx7/NVpGcORhFb03HdbO1rG2uZiWTiXQI
sc47Ee62zvOcIvN/srQM2HdwXLuyZYmwgoUVmTGWMu0LuAEGg/B47DZcEcljZFrw
av/WNBEXNo8gS9FEj9yJw5Lmxbr5ROyLXlvuICqI+5M7GXr4owOApiMhtpaW09x7
Bm4LWUy7UAKFFM9aNj9tXvrfsMDXKxySRAMLXrWLGemlEe9Gc7P+DR73YmMrB+XA
6FchgLwXwW5P/M/YYbsI6Qd8fmREXwo1kNlWqSIwy961HEns/tQZcvA+3z7p94Qf
3+u7bIeA0NPgnj/4NBkZZFvjkQc1bV6qPgQ4ZBgq/i4Uqmb7rIouOZEB6EFZPrLv
4OP9uF3Tx0Vh4txc2j3e78tjwRpMhpMkSAhSot8QzejQoFMVM7gaPRhcDBHMuLdm
NEfF9QrVi7HEcoHewIK9QvmCJmE7Oa6M22Q9Se/63pW0xYBkuoWQCCT90llcyKSi
2RMCk5swb8rxWoPBJwe3dK9rzNL40bh8hwY/uQJLVbkqW/eXudqMSSKbXhZ6APmN
BiDorIWy50pHscyi9UsVZ28u61vpKwMdMF1xOI5yxPyir2I/M0Sg5OnmKQEJoOcZ
kzoVOTyjO1ebe25kqCR4Gl7Ep0lDknRLFv6U4Yj83qcGm2t9Qvs83wtiJQYXm+Ja
EbBJGA0lbwqT2AeqrMgh6AY8dc4kwXu479Y0hs+Kukje1q0lRWrrEaZeZMkNyVeH
AAN1Xb1eWhk9McpDeQ5qTlIkXHE/8NhvDMtvE7UL9XKxI0VE/AZnxm+iAYzx3HEu
9YIs44JGfHA/9x7fEJQIsfuLagu10a7MRBDj59HSZSQMTebCz7c26zn7UU/64/Jp
B0vyw17LqN50abR10mOuxqjDOoWno6KddVBoyJFFq1IdldFvEKCOhQd5ZZbfqzYC
cPva+WMol7izXkKCLhHlH35m+st8jMyC6NhRJQ4IY38JoOD814TLFART5uEUnKnA
LaF+VgyiJmR3/7IPyp+JjYqZ2kpt5dRihi9YS4Pk0BavQKvD6MVrgZtE9izikCD1
2tdcqokKUV3j0/E9PNEuPCYsrDoM6xrfEILAQY/GdSyrO2LdgFGpJpONHhSaGgAF
c2+sFi3HDkqL57sy+7ME39DJc+qzBFfix+gHd/oiESmcyVjdWPiYCp8fDnK9IvsT
IGcqMA4qZy70eIVbdj44sjr2Oh7cBkT8McYiQcg6e5ZcfpkBhtOVyPLmLCcmEMw5
9vR9zTj+DwfoUUOBm8siSX9WqGd+aMI/qK9aBXaU22auEwC238hmxOIOzxzxGTjg
3v/sB8f6EPOwWLuhynQltG1Ro2RosMPdea8vo1fqHEZS23eeObH7bcmqYZrD9GnB
xHD9YfvJBl2Nxvfhv3jmI/eoCD7A0CwxwEfdCajw6zwQaSXydUPokjIcbdKYddJd
FpNuQLv7ruVcq6QIInqBQZFif+5g/ArVX0T4uEYBTEMAjvi02fcah1RgvKtAp+4x
eD3AfmYXIM1F35HTsQQ51QINk7yctADKHqGqnyO8X1VFVZpfIXTrwgSjt4dxH82w
I/X1IE8x2jqSaWAVnLuXJ+4jb1hPm3uyng5hfaujYZ8zZm2GG6EkKqiSaIbMaW8l
G8Jvh7utBn9lswTzwLf0WJUsQotoIkpYI0R3A03hRz0DS9rgD+SRTh3MviZlh53z
jvfEWcIua4igDRl5m1YrBcmsdGNCD+v0RAKudqOc2i7ectAVx56SgLszuP6TsZas
RYKCyUemXaAtafNY3FZEg3Thav4N+YTlYLmTx0lu06PrverQx2gC1qLTKwUomqOT
OsMcbRQ2BU8wuo9wYgx4VIOCkREgge7JLfugOtIyRthf/Nfk95ORz9dllAs5dos6
wywJMZNcu/qFYp+dI/S0eMuT6647CauJT08neqNCIax8gEfg1XT3ZaymSLp390Q7
eFXL4rnG97FGZNgtVmQhKmDIPraCtI0p2aXgZOXM/FUHBJBBHLTgQzPev5VMT+ie
r1NiXdTDHHYeqYj0XubC8rcS7Yxyp/miAuCQ1aGn35KPiZFCloea2y3yX7L37sY5
jU5OvG7Qhn3cd35JcyZtsVuaPSLOXJxpLlQWnEIN7psIKIfC/Yyo0gFailZivvLU
Z9nlR+eEBfoeTy8DpXk94XVZNxD1IikxVm+jQR4SN1kYmj864e+U9kVpYr3OsUcS
potostDmu51O1xrXhTF7CAuj3qp2b0rHLnv/y0deTeVkGO5QMnEHJIhL12HUha00
9VoejuCyTwH/ofphsAsiF9rIq4HudsMpos6bibUeSkIqAb/9jsflZaluQ45cUtTA
Q5vTVWUv/49ggk8/OPjXMihTQJfQKIaMRtw2e2xujl+1rE8EEIm7prVfD0ZskiBT
W91Q3wtVO0Tscz1nLHgZh3vBMalU2fRKsXAYxGH/Q1AbgSiR51EXkvckQaRORz8R
8pUl42xfd3Ch5m0ED03R3oIlgCoueS8sdbi2cYdY0fJXaeQF0F2gQkQW24gV1Bqu
tD9my2pG0gL5bhv7kv48sr4a0kz55yNPTpTk7thyonC28UyQ40sFWEx/9oIRuejn
epdoQSEC6yzFIRE7USeBNHkIYRgeOjLQ4ufnT+RU7oL3/82zCIJKlA55mfelISBh
qdcKOJ8+ltdWdu/UempnMZQwgdFRwATCWb5s4lOspV6IH7q9iGAJz8KFOvsC8VsT
Xqre3aqxDUx22R4eNcW8IAQi3jVIq9pZCpK7x2Zn9E84amH2b7fl4APjjXR5zYPi
z5nZqRhirlTklAkQ1pQMdfhJfBSt7Eb0PK5obb9Hnj8FS/t+EzTIS2N7R+PdghA7
SFja+ceyJcOsKZuc3Sk25crsTBvVX3W8lRVRqIwXTPv7XnSKp0kbs4WVCZWcZgeB
ZgZU+P2mMrbn4DSxWcPzYW5lPAEVIqR4cU7Oy+VVyXNOmF6r38cPC9ad9Ys2Vt8p
YCEvHbx3pniWSoEZ5oy69heNcJwKyC0Zumc+AR+CZkEChHG8RCh5w7o0AabrcTUG
x3eEBtqI6/NC4YUySrdk4x5YouUukrALxVak8BiM6piGoyM95iKPku6RTordefEi
b2PT+tzczPBPzQ0WnQtn2VMfXQN7J3AZI6mvbAvM35A/goYd3rpOFhTMu+9aFrBN
LxQYQXWN4MUgBtotiEj1JQvMnIKvI0pKj+UwSCMmkfDwLTBvoeVCuc1F5OhY4wHw
TAWuFZj3Q7ZTiz1wgSQIq/fRNXqswPJHbBHelLUpcJ0G9FvLXZkbN0kmYUk1nSMw
1HP0fpj0DV6nm1e/ZncSDnfsh46/XmsGzswudhl+eaOyzUx91cl/8KPTeL1/6zV+
8dcONO6s5GvsLZUL2+goHtQjCoo6M054iLv4RiScpIe735kipsO32PRYVXm3BdAi
wUJHmJ1Xv2CEGOcxwXVMh4oYtRcQSgACGKZZxkXjavphgUg+dX2/e+Yw0N4d7XRZ
zfN1OiB9sGncOxzbNSXpr9rR8X3pyYDFBQzRMDdd5AYK+3lydlQ3CczIa9QeycC+
z5RjIxt6sE80WZaaMTTupS7koHO1Eu+9pFShnp9HQ+AczBgT35eVLg2PT1k/lZVS
+VuxJdosGJToU0LlZpiuChgHcsgORVVXC6ugH4fi+tt1aDlTXdXwFW0rXI9FpfKK
GjsA31o8md3dqL5+yGx0nryOEP7LiSPy1gDTnhtpK4XGykGr0V6Uexi4u2N6jhFW
++6fIU8hHpBummtLtJrFcCJN7IuvBE/SUJfpGzdVa7hzGcLqLFrea8xZaD2zLJo2
TplvFfugb0snTYKxPZLL5Rgr7Au3G31KauoTEkETArNapdcuGtkodOodUA0K7dCG
tZXy5kzBAcytwdkzl3MuBBivkW5YiR3yvlzZ4VvsDG1gGDmf62wGjYQmyV0GXkse
roxZKMg6l87volcC3LvJRIvk5/ohIYQ1BgZXHeaRCKYdHzlByFSe9DXEI/oY1vr2
VW7r8WWDyn6WGtXtfqqqovV2EWFI6IfAhbZ4bVcRvKG3w17B68i3keulrtei19qn
BHc6YFTB3v1FQXl5PmestM6PSi3304Jd0RxvJbrIz4UuavfoUkzZ14akc+NKFcbo
/GLIKHBWqMmjlL3gnSsoPtZ/ScxzwsXpuKOdCpLh+kB7enwsr8Hu/D3B3iB88M9M
aq48Wk+k8YNxn/YANtjSGrVGOHNgm5I2Tfcdsv76Ucc2055PfjVxwdHEA0vM5sft
CbRTyXRIB6b0YplrN/cYoAjQDQo9hGg5RoxLO8L34vu9uIsxDiI7ltguuWCnk+pL
fNhAdKuON9/J0oMCkC7aa0KcfXPrirmcUWoFva72r6wNjDxR/hhtOVocIyqMBecA
V15gowI652avtJijhcyZmNWdsUipW91uTEoUQNMk9sBgkbx7oqJGmwY1J3/cFptz
DbIMvzg94GfjXM6Da5TsoRBTwghQgn+VUz+T+iDf6+eNnlMVSBGtR/079byWL+8H
HlbCdSRpjztOiQJCP3zgVU+JyVwngZBRv34gDUqDtVSdcjljkHjqPoCTkKxdbNEz
Lcy9WUxznfeXo7bs8p2z7vuy7ivAie7Ab8qqVH/z/4yCA/fGwcr4fpv6w+F2RYnv
e3D0ngeIPjoLFat8494F+1On4L2o0w6pAr3mMW9Aw6USt4wlFLf25Hop5vt/E7NV
jwwDwAAnBm4QyGHscGUqQUunw0DWtt6gJ7yZ++3c8O5YQJVVXf1IyQ5UdMp5B4T4
dVJD6RFIewDsbfz/zWKY9312mkDvyLzTtjMXhhYvferf2NTUHumF8cnFqUy1mXaZ
sOAWnpAZa18F+JfF4fV0GL2N7rZVbnGVXpesdCY9r/Lmy1ilUVZSpCEqR8uHWK1I
Gbv1B2nzXNPUEZk+NnT6mxzUXTaD/Hp/wya5Q1I4ShHvUA/OKgjvPio5oc3jVo9K
XX2QIWMRMcJCEiLnY0pV645AjnvKJYO+jkQIxgOjgyLzmFEKTbXRGO2DdvrEjbvd
thpRJrCkvUYVidrP7H23AFkBbRMq4RCog/fsPZgDCpW3Gg7iaGhmHYuylBQ/s6WI
LWJETn1kqhG+UhIt8PbfaY4o0cZ00Y+hC4VHD2O+CGZsUPHAXZuPWmoRvRRBpO+B
+QEWO8pcwx90Xle80+pdVmBgEYW+1k8SAasPsNtMBCGNniZD1G7I5bkoi0utuGfs
zMdn3opC0xKq91hCrWJe9udex/4l7qAnl6EWMuagKCU4x48aBYUN8KIYRyan3bwt
aauGezqdFOXtAzMLNs8SPbnu1kVReTcsaepdZaAmF7unwe4zwbtgDbT5DBOxYKbL
bgw1I+y8RV8vs8mc2PL5z3MYew+onRwZIl30GjBfRwXEsytB6Uzt0eoF3xvKwGF9
7MLqnvS+1ECA46aEfcqf+Mne1o0mBy/4fjvmOj9xxU+IM1HcGekK+P3OCgQP519H
BZQ0M0lGb+u7XDhXfP74R0wzWODoLThHkYAkrXubj6SVXW7OYLqYePApst/7Gu1T
IrKNjvI2Ovj8vw+U/M4XDd+aZaQcEuveBJnex0jF6EVD8l3jVBmBuzBD/kB7opbP
XIcutn8MvgcShiyJ59MJWrkoMFOI8L2ypz9EO3KFUxUDj/47Pyr5vkLvlyVo4+82
btSF/XCUmk5ZH9urPNuhptPcXiGMDRsxLvH4SrkD2REsJDVX2qOhLQS+LzTOH4GN
qiMKpWRs09Lo8/MxRy5WZPD9GJZG6m1UmOSJr8xuNyeIFpUtP6284qurcEzT3jlc
R3mC+ILAZjT9XEh7Fk6aHulF86MzHkwN8uQSi5MbM8HwJwxUjCeBlGWlW9pweqQL
xcDmEV/c25MU3zfIEzdFNUngVTmbCZiB7CSUBRXgYoiFFVuoReGGeeye3ISt7nVv
rBpE0+BCkslNIhDYCrZPm/nctIPgmFx08DMaMryavyRYMu943KSFx//kc3yWxW4U
VWQiKLeAAAcxRgraTio/XtcseBd3NNUD8bucOg/kib313oTwJNvoGV+plL1q7PiI
e1bTfsiQSsXXMHii0GqE4Tt0xmUSV6jaaQU5oSDdfnITnruqd6HPpA1dPfFyQTDk
hnI3oCIKqw+slSCjmIQuFVXnEtMxN9sHZWHUb1T1ToSjPrVe5ngeptnGrwzMEMr7
X1NvHX8ZX1pAj6BmNFiy12xPc4swrB4exeV7t09FUWWRuw9fJ76c217W0LDcvEaU
lwnKjdqEP+k9ILjR/sb2C1Affyy130/HJUZyA1+gCPDXYkV/Au8aX6Q4rf5ZmIJA
HA64dweeLGwt2reeMkUVeuSdQCNGZWStmcnXMCdxFbbbigpoDwd/xfSK5EfluCyh
YNPDEyuuAYsyixHYfjkujxqowjVgzeGTZbA4Jk3cV5YYArtEUcQxKc+SOP6sez5V
Lq3J5g5KXp57XlCaIU7idulNu+qzjZFBuUidkBWLITphxNX1tUFx318ujr345UYy
8IoQycA/LWXlaFrN1cRs1MULNCAFll2L9dPykGPNqZHXvy+e4CghJta+rk497n75
swwUtVpKcVwcOvIOQKrXdKB3MbWNN85fJ0MWuQIoEY9eaQ5wzidyF7ocAllc1EFx
+INFjg48F11c8a6hmC+zC2wO+St26ed3fTa5J5VigO3/glNyezZi3qiKnWF3pBoU
H/hvrgrz6l5iKhZ1oksFgSs15cjFdiMvYh/OjsQ97QjhLWxjifOy80U2xiH5Ifek
fjWiqPD6PLYrGAPN26hIf16mLxFYUZCIexvKAQqXHmNPQGiiBYVOFgPCutqj1ezH
VZPT5uTzXUJUqAFszMY31KZwWtMbYeIB/6UgxGK8OnMm+eM8/nbk30jEuewocXYa
L0CMK1WhEPI3nLrpBkoZM1q0xPs8Sb8VlAkXWAkZ+7X14pg+EcC6zFTYGAb+WCjl
E1rea+wawYSYrxrwSKfDaFzXtvWSH77G/c2VPC2+xV5K+pBBHljCB5GMJzFQwbic
t5wtyAWKvks0ouIUAQiWpro1sbose1latdoLl3PhBURzFPfM+aZPWSR3l5j2wX+y
qZ3l6YnoD6aTvM1Bl0AIMlnLMXpFK/+CjK4mgdWw4SI36xq9e6lnYmvg1nFZYvZp
qoiOlh4SRSPXCq0I6CEX8zgHwAcc4ETJ6ai8NlBYi/DW3GFBFcD90XC/j8BKG9QK
Qs5XHy8huS7RyEUHuFHQnm2yDK68ItpzQzimDULV4aodq2aORUUBNUOcOXqLenB+
rHtPc+FQ5Cm5aDHvUWn9YEBXwP57jV7+vMaGjVlqQEjdMvyMfcC0jm3ByKOUAigi
hfSHTaAEk31GEuxjtmDZYYFukQZAzIXoylFMZtZ4k/SrQwuQIQ4aim2kv+RRdePR
0XDiEooLf1KxagizFNncXxyp0wQZFvEXdMQzOZgbvxyz1Pp7O9hxHwtsP8aSyyae
QaQub6+uxwu7sKAx9fXb0wv23J0Hhi2ZLI7PKGhBgdSGd0/uMz8ocaAWER5QcLP1
o14tAFei0KpTMzp262Fe5DvU2zW7pVLFS3jSgvnY1kEKdUQnR5HLRBy3ipoWsQny
WAD5qSSWO/M/iAvxNdh5S++Ba3cQ/h5yPBTvVHOQXi7wnk8Rt5czTj/R8uuCuNVV
I5R6Jo7oJuhXny0xvUBlmS+qYiLOF3AFz/3nR7BU3NOUPLnQZTtlZWgK39B9qwMW
IdjOyGJq1fcEk8k3W+z06NPooZsEx5QvwYSu47G29DwHH5yptS0ZnUGcjVhHaITt
6V2jnF31m5UToaiuvjnTOxlqDcADOZ0MWZOKgM2AUS0qXnupgR5kfw6sVp7aorp7
qE4ZJz90gw2wdcYjrgJTcVOU2tRyX7ivH/TIqIjTqzXyUyoMLh7GpF5esDdHeZBe
ektRGEocZFFVU4/hczffLcfUvs67fBBBnAdMcC8mi3+HqB5Kul4wZkVIlXkAHLri
HSBA5PYNjSVk28pUQGwRyKYxkZDa9oxfX0MnSv/62vsxzrSoctjR+o3uR31Yvmjh
XtVEJqxVILDDMKqV+w0k4ZZ6REFS5ymlcpOZW0tnrRvV10v8O6Aapw8XilgIMn8r
TQA+dWivL0yz1JpgM2JDDstAmtvpJKbMWMreTh7v1bp9khDiz0trFK6bz2SqAb69
bE7V6faYxT4ggijgvD3QZ7VSXunAgMmE5NGRQhFZHeidy+hkg9YBML+t7lwWqr7T
dZ9JK8s6IfI1RudXKf4P9XJCpf/eAqH1bJDRJyrf48yDun+14vkNToR1k1hljgyV
zL9pBoxJacGlmLrQKo14jGVMo6odKuVTEmurJAoUk3QqIk6C+L7DF46sL5beUTWG
z7Dp7HgOb2g1sXhYfxYbwYZnjYzkvH2jdR3B04EQ3tTiChS8Q3BVssYmFuQiGEvU
IgpPet8UrliUoUMF1f4Xf6wMPFVbKIrGu8jXofW+PV8LUxL0EJJ0GOPhCcE5a1C8
eejt1xGLG5Hj17kTD2NeT2viVmRXkSaHYdAMFnySV+GY3Y4YF3yGZs3yvSnehOxz
6JCDqL7Hcvgfgtb8UiO4tEUvkZ+SKa4Zl2i7OJzgvozwuDzwXFmvQhZCeIeRDrpV
gaKoJboZW68bfimjOzrNa5qAc7bajvcjgV43kqYe3WTcysnWey4S2tErv04s4/kA
y7hplegwb/dQlKMRUNcx1soqo8Kk3b2g8CrQXqG8j9XlKVjrGRRaywTiO5u4oT5G
C3afLzV3kwAyNUf4hXXU2kqv73DRJXXLx9rOLLy9wxAw9p4GFP0glwDLBMZCtE8k
vb6o6kh+1cVe+uU98hVyxlNIJOrIHuJTAFvXk1ssWVZ/C/D3/QFdWtDYNFjnksFP
O9YD+pI+rCy1yDS5ZGg4CGlTInjF3s8x9eUHbJ7ee5xRGmcZgdMkdu9WaSnl5xbA
f0tBfioQugK9sMIuD/1nIG27Oi9YfhG46N9jbfG0fGHtC7rwu+vZgZxqJe+6phcE
rq0M+al0CC/XKYJhqtNRV3gVwMb6J/Wr2JPhqlXrBECYZ+oabNX21MM7TEUCsYRS
kU4tuBaiyEDs5BA66XpuKkxtxlcXLj64ad3E7MNSuxlkuvfECJneM3mRurdWruxQ
l04FPrwF6kAUwQLpvgwxwdAeGTr6mXlz/bInUcyEBHWpUsntifcguMgEV+KI0g2I
n/f2/a8NxFOx143yttdjnUxSl3HlLrbqZp+Sv7G+TUVAmgdFe6aSm4i+Q7h/ZvwO
c+7na4IZKFKLKo9X+/7WY6f+Cn5+YkInjv3iTkXG8TpHwNRX0Kh5loIb9E6Bgwms
6BrUr1OekvpQKgQWzFgs7bsVW2fs+qw5t+XglwBDw247Jt02RZKgwia+eKWfG9Py
SlUFHYDDmxilIdrgQ5ZGAbFSgqCQK2/iY1p6TBw23XpvfTyxOh4cndDo1GXKfVMN
rfIWZoORoCMXEv0GEhF6q6Yk2MSnRI8bvHcFy+HiPfGNhuQcygPhLLNkT9HBNTes
/ubSg6uokGdkR2u8X76eOqpCxPNRsrx2VAHwr8sD7OkrH8bBwu+vpG7hGOnl/ZAH
Ni6vW91TQMUeHVFg8g59/B0Lee2nQE0FRLlcLk76Cib456hvrOS/e/hniEBWYtoU
6MLDzNGiryVIW3duVlUtKjEZh1lmDiMR2MaL0rmOopG4otNuwosKYL4bPgJYQBdy
ZcKPF5x8MG0tTv2IL6yY3Y4gF1QLln5/oX/18flbr4WGk7OoXPLqY+402flFu9Vb
ZOw5h5UvhLxFYAhL7olWoIFJbR1PwuhPEHwHRJdo/+4AYjbUEVQa5OkKkRv7e9VD
CHDJNZTwambiqYCL6/JDeqcC/+V/f/wSIW+YqMLejbpvjyIGm/qeT9pwOG2KqaYJ
mzfAN/DoQu63TtIAeFIHnvE5dhnDLguFCS1Wm1lsi73zcaFYDRoqDGelfjwzmgn+
WPBloDHMkSRahJYPV6nUJgYs4W7owwZ47rpA1fZRY0PcZUkzeOVjxAvnIZzO9Yc8
1qESESnNNMIzeqqXRjH+1Nj1dCDgIjMVXWFVtdBjjKCZomSNx6LfYrZMQGGAI+Pa
dFSPuSED4UpUoRGApr0ZIbtjaEhIieSSkZK/EQROqXSnNYX6SU7QMJHHBx6iYqe8
DOA9t9zE22uO2VDEo44xehf3G2i9Bx9D9AbSpdPkKE5xQxWeL1WF6cFsClt4C+Pv
QB17XL70MN24jEs4ugNprD2QJQLlhtbunFnAN5l9TwxB2t6elpJUy5Z16ndr4Ds5
IblcDcWy6u+VlAE6iLoTIsqL5q02sS1RivGMU7DF/3RqCQUO4HgdQs7Pr+FTTs9t
X/1FqtvkwJG+FqMdXS7cdZ1WQu+M2K8S29DQ3D8mYAFv+9qOEZaNoYH8oF5Nv6jF
9a504S6lWdAeEw16/wa8o3bKaQPKj96/bEtBu7lIlWS0z0kBcc3uVEHj0cLkrHx+
6rAGJNpFrf6fzAEBBYcSDdD0E3Sb6/aYeOfnaYOUMRr1YK9LDXeNT8FrsE6hryI7
G20+fxIj4zkW8Em8ODaJZhZTSGAKyRXwmVoHVln+BI2sVeDQPZQ4rUihO5gteZVi
hopaMf9nA4CBPOEYJ33SW3jOtQcHduW9cI6IGnIwS6xs/0IphHRICQMKN13Rs/G4
DkiXUiDTaBECsmN/soqPJWajzSxofWhLPzaBtt2BW+CDmM/XFiYUcRPWbAoLn09q
6daQJPIFrnZr752oJI0SNI9FyDOMsKAVyRACg94yYNQb3l/6UMrN4cD17O9ARSE8
TY0c0ivz3El7H6zDBkQMjfBOnzk8EqMRzWr+5sYjusg7MdsQMF0t1izJdlNgkLYj
qtr9HJ+OxHY3MucSQknr9DL2M/65Ved648DrSYR6s67SJmVM6uTuEEKsdfWXjFOT
ij6TUJ5JR6TUoGCUvG5aB+nudbWYhTcD3vUcGfYn7KiZHbHVdI0VxWGm17995P2F
bQDRyBHufNlIhOVSqYy9qTlUvxgGlG1WvHWytK3mUc1LvA4enZ8bAppvmoMtcO1N
NpYMtUkNsmhsQoNQDVoz+PywrhLAb+ymyPp1l+nxwk2KVNsI9W+X2E6DQtn1L26W
3v5t2PiegEb6iGiWDD08z7z1gypKBHOM09TSaZRlyub/pjXGrgNAUn7S3xTQn/oP
7iEDZhTqxjw/BUd1eV0rMeQylNHGPhytFx6d+q0i88QNT+TaqrSkBFeuLEU265oz
FSh2Y9uHHIVGglyeeB8HysWEoT1/08uq4pgmfalrLJZkR4Pn+uytv2oVdkzE++eK
e8xqWi4jRPGdFm/ATN8wbCIZMvwk+sc+6WMxHBafXGMxyKdPpBSok060Zaipklv7
MrkLf8UXrqdf/lKNTfzGQOjwph6ADdtCb9mPKgDapUUk3s4FG111gjObIlkCFTDp
jeRSpoB6mGIKhnco7Sw0KnysQzAYvr+S4qpRikj1jUrTbijzfPdut4bvspNDy6s2
mVSt/NvqlVzc7i5chhE2rjCz2RWLOqFWptdDJqX1xbBCCrdXzop0jlLSATGSz9FI
uKdN+ekM5+GjrxOvoR8CWUbSzhS1dDI6bjt2WkXAFbUJfsYD0PQJ/jGlJjDsPluP
th0yaQegfONL5lb7kcadusdN5eyCwAAcceQ0Nt4IUnnzGuCGLb9AOZDLWoTB4cCq
LUN/TYkd7ZpQOoWM/zHIB1qm2wNi2NxfirIxXMAP8QrUMer9PywizNcAw5QI1MZj
mULO8PzK7xBP/DI034TB3bz2UNcyNHQKyUrPoNAFKk26JDWSUR+tSpKYdwmb2FcG
B7enJlzhZZirDmHGO+719n60dGRrYa0uxnfeRcDIVPtVFnaGpystVqtt91DWKsGI
CYVfUVlwZbcqLbNEDyZB2mlDC5S+pRYcMxYR0EAjwEOMuOJ+v/kcG1so2cvXrxoO
0ocP4zIo6/bzW36A38PIJUT0zb4ZS0C+g5+eUVae8N7BUoGi5gnSZdhRGW8/MqC7
6jjc2mprHv0uJcFdV2ZSoo7rBV7sTzQvPT/4APFXkkMzx/I05qn4qPSm1Sluv5O5
B7Tx+Sltd9fprZe6ThPrGoW/qSOe1IlUvl5QaqVvgloKtscQKy8GicMVulzmfgPR
h7WMpCL5QQIP1yzJlbNyy5fWbD1aeqlDuhcIZeuXvzuFsBMJGQbudTYG45c2X0p4
t13fDn0wRpGNPc7SjgpDtNHss6L/rtHEaPh2u+FtoTRnR5wORzXdEGEWDnSE4iRa
C3FSatwk0k2WzU9S/bWGpFV7spB7aG92M4wBNR5MP6GjPIG5skFHkSN7X1PWEzan
zdGBezWveOGl98hhmnP0pwv8Hv3JtnXGd/W+JvZGopoMX1qH9Zlh5/zlD2o60KJa
tt3SQjh6lt8DoaWVpbJSXT1NLA2zFAMNDxKjvl9hqnPG3gvsQ96ibPwcABeJdjnw
A4hsBYYlSGZv4qKKYurDgiqH22vhrTWvml8DGxdy0Gb/wfz9pR3ODqWXx8rnyNp+
Mk38QWdlcvYek0dCSUJ8IraElm/qcdTkuqKIGT8mRFL5u2fko8ocEVDlabEqFePm
TY33VBA/niUqvyQHMGx24MfiOAcNR+wi3pxev82FEGaQs0IYBhdD/bqj3cMoeT/5
gUMuHIUp/JYGOJZprsy/zUnAkRBiEMV7L+laEg37p071sESLIUnG/m6qnU3tAieN
qKK6KJqBZCv2tmi3UESuXk29Dv8EdI2g9Q1YnzNSc1vxjHmOktp6c/JhwVpQOyzW
T6dTskW94saxpt82NpRMLVFojp7vjOZOG3I5miMu8PXyhZBVUJtrF0JhHnon4DE7
J2qJ91wJHdVR0dNYIbEMVXbFHzskOfPDZxNOWoP25epPKPBM9JQ0dntY8gJA3m5a
hOkfzb4Ea5NvA41krdyFcREwtKtI4W1EvfLG8am24yUiKDwD/LJ/WWqnUNaPwiAm
qClW9MYEYBCz3kKKOXndKxFFot8CTpznek8dR7yHPAp0Oh0YgNdz1uoDR1hQrvGM
khpHFm4gd1yuOQyn/SBMCVaJGwDRGACdcOw6d6t1iNP8voU4rF1IFphphFoLlL2n
rDBpmyIzvCXH5pvza9offEICJAe4HzId1EEiSCE+rGEE0W6uFeuLCFv3KrcK5bqU
ge05kfLECm+y66wazs6gIcaD82wGDRvfwJ4uL4zjC4kNs7G5uFNdJtChQUb0ezDx
XKoFuyTbYdsQNCntZn0LnRm4MnIKsrDr03qDDTjnRaTZLczWRCJVkt1L04dB2Hx3
sRBruqbrXxL6ckFvSJ8pR/2PP4jU93HhJpBFdjXdxyf5fMqx6SxLoKvypaGz0fT6
D8GwR9BgQkmmX0dT9acfSnmeH200/n0gKB7wt+bX4uqGNsBcQ58/pO55ANXqrAze
jkExO8Jb/UXc6CFMOgjgvgXbYohKUcJpXeWiTvLsj0r+LnSZue7P/F3fqmOIbXAq
v8k81gNgTT0GAUCfmSu+opBk/FSL6KQtv5dLlNNz9MGpdN6IFZaRcVYIA90a0LWp
ngQI49/5jb+wyqeM2ghoVqipvF6xRcXN1y6rnACeJKodvjHVK8IAFbHhYgFWp/82
uOw2UVtlnI0V++NykSWM+Rw61fiumSmq3ff26Q2GLAcuYNBdGz26vOFQ1dyLEkfm
0LcF+txofDz0FBeWjBqR19eI5Y8VTK1qCQXSrOD3OKZo8qWpUpeWQ+sVnZexpnt4
bfyv888YBLMY9wuH3ZZmCQlaBPs6TJFcqE9AMaCE6nQvzcaDklUxG2G1eXhWDzQE
JBrJoxhcWz8YtkwEzhQcGnDrwtsro735Mbed1hl07Y5nn6F7uT4K9tdK6PJJ7kWo
4+/VuS609JjMtzqvCOKgcSUzC1KPwBSn/dFonta0ZaI/62kllZhqjGwT2Wr6Pf5s
eezAdlvYezHatd4ZhO14itMxAdVotzqJeUkc8HD5WjT43Vo/Tln0PuNUwOqICDq8
cPJ9fdKQOTlFiY2zAq/94sU5BUoL6+LxJqsZQQ4KgcLsXHObtfChrZBuVE94y9cf
CD7BTz+S0Nbe6ICLzDptnxBlFQws1aEXsSCZs1Hv+MKS8zDb40WK9S1Kjl6MuboH
ou33e8BHT/ZEp67djEmrVMABEyKSrvRsu6dIXSJQ5jfCw6mKn4ikID6YDLt21I/D
bMrJ1rxc+fJo7CYY9uapmpg9VqVOV+U41erSUsyxu5O0XSmBtix3JGvoP0OaqJWZ
Z+TtVIRa959uhv1iFNxT3d+YXd7JN7QpQeLfbWk7Kkz3W4ahJqMkfhnn1zXkCd5h
4krDHQynCukdq8rOj5MNOBAZANr9jFntqoxkQoifRasvEtPuX4+dPzMOCwuKRrNA
Yd0iCRibE8fVsTvb2FwcD9aCP67IVWjMPNLm2Umj59k8m7vfn6+Dceg18ldRBktR
zt+etzQqLgLIW2V31QwBQJ13Jtf1HZtZ0B1Db7NFA5ysWt5lf/beDngED08a1S3L
qJeFpMsTP/WjUOHoqszzXmlwaI1+MrJTTo2lQx7R+Xz3ee9ok3NaF8dbHXfpvGPb
qtyDc8twGmX4DSnvTDeFioDUGYYHWUK1REQslI0rYzYYhs4+Dob9IScNeF+R72iW
dhuIv5fe8X7CTSxdgro0EJ8E6pu4cZYLzxRVrMppDz+xGRxHfv9Wwir3xHBd8Mai
monhM10mZSWVfEXcKoyCSaMYmmHF7RKStYUZmcXpdYr8nwquR9PPjPfTznUWBQTL
+n05dlf0nbqKVKX542x3zykGbJZ62V8DRVj3BkTjoahBeco8aGl1IchqdxVsFpFg
Kx26qu6mB2XA3qQ2RW+y0EYAE15AdJpFWeiKZ94nMgjUi3zmkaRkZw/poD8BeGZ4
ZyhQPEYj0/0DgUdHjSGgm/HF7I3z4coZDbRRIOBS1dZnMBpVai630E5pha/cvjEK
Lq4YlAwi25vwyvYBJXfMXqqGnKhAy5WAwXbALWqXhVxxT8RyJgygyj+vbAQ1s6G2
tbKgF2nKwDdm89Oh0XKofBS+hwMIBWhrZyqgHHR1xN1/UsVTgyoR4avuwxJ/miJh
5rnXWbWEb3OK+pnCIn4UNsJ7HwPvLPWwYPrH++0GOOMaLXe5om3WX4IQVtAAgJUk
m2U2xtPuGQCiSvxRlj5n7XXD8yyx4prS61u2BUcr/ve/++DYI0dvPunaJVOkzKpT
xAfXr0nlBrEY4lX/x4tjK8uOFsMDJ68dRUiIJZHXntiqx1snlqQVEo5r0JtXF9/W
jvOV17gtFdSXCC6P4hy8MqNNrRmsaCbe5BvmpNPInJgr53a3+HbQvZp7MvjmGSwQ
OBnbbYL38ju4A6QqC0IUrmxnqttyAXaPtWuDwX5uhlu+o0gmXFOkJEQXHBoOHDHF
FT6mwV20pbtpYggXlp9mM83/3DWhEvGexd2kjFINR8tgPojb5f4NnQ+C/u+u3YRC
UJMFJ1tqURXO/POt8qLPxqLDcNdXmAfYrZBVgqBYuef/FfS3/iW10F2ocHoJ0nfv
86g9FolmLS3fqwtWGOxV7MnXjTkFirqV4PTN7Er+Abo8ayNKmdPmIhrZWs4VGeqP
wQQzPzBrmXlSvp9hmO+oaYM2mvXnrPjGDndrj2koJZVpnTtCY1LDxWMpbusKnH6B
bwRZ3U9iCrTUhILdaNFPIy85QfAyN5Ku9ECK/Kf97Q1RTay/y+fgaVXfzSQp6j0M
h++mL3+K3FLOgT8Olc+JtnCzCt2TR5q14mEh1lOWon2mbrrCopm7aa4vz5CDXCUZ
aZsrX20suZUcL0fPZ7uSlZ0NRy0yC20N15e8YRP90kPnJYlVCdFBoDASOpJyUxDh
LdwmaxwkTu/AdtZPLHWfJCZwwNkWw/ixQor37UB2Fx1f8Q5IOEtuS0itxJlaV//h
tT1XVKaf6H5tcaRBhrITL6NxiHPgJ/EF9ql0n9Jius8N29YSkDp+HFzz6qtw7Mz/
AE+SoV0o7p8EJw5CpbU1/3RI+b7tzGy/Q0ikrzJrK+LiVm+z4LXr57jOxNw5cIrI
34asHfA6dnHp7sKfWiQokb2HcIMwZoLHj3NVuAwPiWJsrlygt7vT7953g5B5LnYG
vpJXXHqUVmA5uGvJt/EqQwp2Y8kaQpJ7bK9kU2A1K6mMwdTTPbdlVcKhnRxVu0WC
NjYkoqbX6J8f+GYJ4LW+2mY8QaMnzQgaOiSJzRG5wlBPsPZ8xJvh/LC+oAIyUlIQ
pGg0LqYng3Jbat6l33c+4+gvNp08Ws/Wm5PML5UBEBohO6BDQHA+UccJsk/3MlnI
YZ44uNZCPdhBFJoQHrDEKp7ewAkqu2I4QXdsEWKzSF9yx2uJyqRwzkdUqMilLd+m
2gl+PsNzJJX/kCskk64j4VwMZVuTN6U05rYAhevZhu5ejPmENPdPcR8/S5mlkMUk
inCdl0JBtVHU0nR5Q69SvKEy1oqGf8pIQD84chy53kJbvvpY/9mrwG9UxS6LzsRQ
dq5rXuSqhntoRTx5L3xDFSbfteGZyl6KZcksN64GlIt/fwU6280SkemAhz5+6b5R
KQShxNl5sOKLURtbUPanFTZdm5i+1IrInTMt+vb6+imthY2RinnMIsShnJWrQ1BN
k5sEMsQQXtLgyxLMmI0my6//GKBNazY5Y+ugTKTaGS6l3yME+b9AWluGNCVl4eWm
ZlNEYd/na5P7gaW4rMQxBtPxtlOKt41sOEFci9kaimugwn0YJF6pM7oh5Fmre/Ya
WhA5AukG3zbFplrcU2IvjI2NQUNovIySRxw8fzj24pNPUMgMVRUi4T7iBCFX7JQL
ea4sMIXV25lBFru+VSpYxpntEIgsrLN582soaAn46sHaBiK9q/TAXkHwYVu7CE5P
NSNfsrD9FOjuu1TVjOOQxI4Z/E14Qe97UObAP/H3qVeebCrIBzvKJlO7A/oIw/uu
7fKrEl+JflzVI0UIUU3MH4hiAu49xshnCscUl4GHurZ/TA5f33YRdUHjykDL6oXT
JctV7b3mqrbC4Xh++Q/jKohQEYhCEe1UU5dvYTVJpYrJ+GKOfz3k8PazxGzCAS5r
rZYX7Wgr9uBpDY40H0Tc6Synjmx+p1SEHI9Tt88BLdaqPcimiAYsMVogrlhf6AIa
IhLT0GukF6OUXPGXJlYmSRC36c/YEmcFv6FEmT6mHNPGIP3ZEl3s9OdpTrxn4GtA
eCXoGLgRO/wLkS82hkfOQp6RcMR8DGFZRH/DZPu9NZOqnDDhGCsAYl4m7ZRQLrAn
dTvjKGSQKA2fjsjNE+pHr9cCI5U7UPr/CZa6JNjicFeDU0kb+wOo/rjoj6B9+B4y
8Tm/Y6G6fJfziU7EYMKztwkQKEYUizMq28ta0Pkbg7CzTtwZWheWmzXUyWp7HS7O
cWuEuQcm5gnBPpX5uqJFBQfkkL64WUeaAtKCjAbOOg+hwfqeh2VbMLQkuDLB2l+h
VrXh39KfkcYI9nUDcaSC+azqMSCk62axt2hRlThJHkmoqb7aZ+RIohW9SjLeMEpW
moFjEWXYry667km2sZWkJzbSgz+OCtxW1QcGc+3aM/vKe0rH+6knMfYzjPJ6NhiX
Ehf2e7xK7G5cV3oWBCPUgnCu+E/4vsnZ8OSffCf+vDAjsa0y9IZNT9wJ9xH+XJ0A
//251Z6FksR8C3006a+H3XZ/5SMae37lVnTXasZ567eezEgmO4k3ctoFo5zq+6KT
Yt9v0s7y4tkReCzc82aZrSpxkuMC9edqhpkDjK8Crd4G5u5esV7fkuLBPY5Yv49r
vlzc1J0GGO3QlL0qFUlueQTplq9tzYS/UzNmX+r9CUFWg083YxbClZ1OVK6Qyx7S
+Q/kVZlOXYa6OvBg71dieQhBiE+wbfCAJvA5IcxwZS9zaIgKaZgNPudqh9ywY9Zs
bqggYhIlFFFkd0FSfFhsz43xLD+YIS515G4I0fZKBlm4q6Wm1xor8sNe4o177XE1
Y8ayPFwN+k0kD8CpApHI3HrzNUW5jTOolYzw9Yar1/vHe/aAWQIihsTzSLHQG/+Z
8AVBFUD9IZynf/qsg8z24BABfTgclpeNlwm8L/c2Pw/8kfq1MOA9C21FOb561FRW
HCDp7yTQ8IZxd9m05rnj5Gqh/eiAQ0UjcazGhD0DUbY8oiuV/MlhoFUrfduAPHYQ
ZOkIq0vc+dOmxs3YClX8JCkxT8Bdx/k28UldPEBRq5NAdLqhzp/kJVIaB7vnLxhg
knGV7jVVbohd4uuCqC0qfOHje2TgfehZ1hGdvYBNvcjnwt5zNr/sWYzSdeQna/76
jxm5ifF4N8YhrN3+zU/Qx1yXgC9/0wWGsPY8CnWZY+fbwZYldZUXe33MA8eN+gOJ
fv4BYVmf0AcD1vEzS+wW87ZUKJ1Qt0ZOA6+8oBCQk5lU+bnSZnNMF1cGLSPN9eWt
y49iiOBBaD6Bw/2K0TA1gqSMvcsA3KUC5HGXj9spzMlsN9SVVZzUFTRu/1AUb/SE
9cdyNJeDy7TQseRfAmiehFC7qBPedrKsrRfkMhxgKlzH8Hdxuoyemiga2jS6OJ5b
e7Qly5mxotRMMJtkMN/JmAIwoTk1Y7VpEHeO645IjFF1ZzfJdIYh7+yxEaVz5Qvf
rk3RV8jlo3uwkPy6InGL9ohmKQae9oRtpiYSJG19YlsUXnCxLgGEUWfTY/Mh961n
CBf8wScZuB420gz0IfYygG1mi8zT3cfTgk6mbdo26fb+ZywbCDMdyBClYaPZzHKv
DymvOdPK61/XWNxysCV05Rq7gXRnPcGUD72dJGYY3mtGqHUinSrsvX9pHnDv28YF
aCG+bvh7ipVuh5FpD++l02EMW95h6Ug4GknIx2NAaY9YOXdFe0cyqa3/psoTPbIv
ygF3ItF//GDQlrciDGDe0DHPhQ2jZ+LzB2jRv+te734QMw8WLR2hfJCjx1z5VAoK
zxE0tPLoU+kaGE0bWsOTiDpZdunOH87MSycRJdmnW5Y40MVGCqrhu9ogYw6dRlNI
QDUo7e4qhREEsLlMT4IUiukTQ5X3s6F+64WC8nhIfc6s0SLy4gkE7XjhH6DsFEH3
EkEJONKavliJJd8J5LuPtGacGxYg+LlMjmjXzdoq+sBAMD59VlxqbavZO9djzIYf
EUnE5q3Q0XLe4FzT307o18HTovgTlQM9FRm7Q6xHXEvYFt5j+WGBIhFX16we7hBZ
y+PrymgF4mskjaW9IIxVKS0lS15jMhduKcvRv42k0ZfcRG3UD3/F9Oi0Gwdkgxe+
nY5kyUJiiT6dtDwocUAc8dohIsYk9tCpAhah/arafjpNa31RjPBKTOhypM1Z63a0
kSEfndNRpBzaUR+lHQn+i5TV793AdzGMVyHxP+CznBN+iFFIw5GyxYG0Sx/pYD4y
8D4e4ARfDXLyXYt1+GANw1gZJpIud2vebbxrmto1dvK//7rBrTjLGWqvaEmvbL6B
3DxjMhpP3UmHK+id5pqSyZ5OqAqJ+PNQDgcsZiunOuv2+ndIMc4l6cFUUH+FCYnS
Vs/ZreI76ULLKhXrzMudVr+uoNXDqL7Eb0r0FEfHHTpsV9nO7XY0XXthUUhs4qbT
ViBA1d0eQZe+eqWxZdcRqw4jutAPbbtunUeI6DGMeAtrbNQ3WLjrZc9V8O6FajLu
N6AQiMzFMW5p1u6ZZHhokX8qLRhUk6xmbV2Jt3GiJ+qIscSZxB9JefWtctiJx2Fp
4fLo8VaRjP0YUyVRt/3KymwMnErMkvo2d6nQHkqzujQ9qhoq5ICI6FexZgoY4vvy
wNhxubhToJi9hQL1BPDm04bO2NdHwj8XqU3LauXG2CG1MMpuIGjcKz2DKAuZ84no
9Okh/6jb74+9Q9alVhocbcTNmmitSOj1eD2bP2a1p2PG+lwdj08/13NLzZF+Sy1L
DqKhRTqsvovKcBXM/Uka2qcP0aZ19uXVr8RWiVAOU+RnELwIj+q4voJCWWv4XiZI
Q2zL7lqWEjH4v8Q0J3KCVpGb9UcI8oQ0cJ4N/hPhdgZMSRCEJQs2USK4+42qoZgO
B96B4mbKW61PSNVHEyIlGy9spwB6132WdIGViXqDnk4bmZyveWf3g/+vHgxIdEg1
Nsvt5I+hwrv2mPQmIhUDQcw+3u4pKwAIPUQlHICox7+JUmEmzwXjXGQC58xasB5u
3XfKR7dBz8tMUnn5OMs272U9kYmJ5LJXT9Ezqca+Cw1aLnde1cc9fbHK6UofDbbQ
vzSmhgCCUZutqmbs/6J4WU+gVcIPKI02ftKkNtpl/Ovipf2QtYPk6c1TKd516uWX
MmHXRDJXA30g83RdcGC/FyfAZlyqtYZpaX4Uh98SRg5vOCt8uo/pgv2S6AcPNBLD
ig2w+HFaN0gpfG189eHUOuf5IM8rGf7kJRv9v61JVLMIhbt8dJcC3cWbfcapNxBZ
dLzSmHUwQB8Y4YLCQ11SBreCMeVuMUGvx9f5Kr3XHyzYNoDdBCYJUIsViZgZwMXj
795zrdvbIUcm4zsF6+tV3MatqSD+GaML5c60SipT4wOCGsXYJrbWrXm/nxLg6V9T
TpGrQF5PVlXMBR0SFPH/zQZEvmMXixHpCX8YrOmpYhvJm3Y+gFkrV4lv8CKGdbPG
liHp2xNMo/P+dRHMXxCtImAzjGDwx/V66Z9We3JrooduaEQycg51DQEBCQoic8G7
gIFXgD8cHPbS7WXF5BSzjJwlEzAdFDzboM7v0dlOGLd/k52COGtp72DgfsUws7fb
ucxQfzpsvHnqKg7Ei83pInxbZp+pRiWkdpMscFSq4z86RI79ZHw9eVL2DXYvmS/w
0rn6CGA5Mkq0E5vop/5gfZQ7IF16NS2a5P1XmnjGlln1pamz7Z4AxDOo0OMitBtA
iRUnB1bqfGt+KLjrZf8Eu1TKDqi+/a2Jbd39jBo0OjcRVOwT4SMEMyCrsyegSGma
9m57VzqHqBSg+ldXwYhLL7HBbSsqHQDWsMn/yjDh2hgRMmf4NzIxKWA9thb9iuZH
dX11GbmZUgsdkbQKwU6IBvJo8gvw+sp0MHRKXGNkethcOXMCDaAJi42QhcLlig18
MNj8UQhhgzksKNNJnRbh76vi6fMNzmfdRj46OpL5IQ9fBQUI7j8ag0c0m1wZICdq
bxusB8Z7s72eNzbNx4Q+w+vF8CsmXpotAtlIs3LKQEvckjDrjP/9WFCRHLKck274
SmZJTpgASL9qqVz9iJytUAf4h67GqWadw8rxICRWUuFtkWIX1nVsU58ZIwNjasuq
5UyrLPKPULa3x9+u+zvFECz+YxVVlOd+ILYJrDPSCWNlJYndoL7Sqoae16zPF0Xq
3YPuuPjJO5qfe0Jt1WLVlW/8rvjnbWdOvVWkeLT4YM09o7kHP903u8KLx7sD+vnp
RjOWO3k4RVNUPRzqjdBJzaGrqbRubYqDr4aHv3Mxf0dACNNmEpcXGtQiXDX/XwOZ
a50At3DQF91Xzt0itEaTUdjEHoMd0EYS2gQQ1u0wwU7oW9w+LLcimw5MoWGN78M4
/idjPLzwH2JWMr2esBW1hh5GE71aKRwyZ2pDQvz+5ag=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
module `IP_MODULE_NAME(efx_csi2_tx_top) #(
    parameter HS_DATA_WIDTH = 16,
    parameter tINIT_NS = 10000,
    parameter tINIT_SKEWCAL_NS = 100000,
	parameter CLOCK_FREQ_MHZ = 100,
    parameter DPHY_CLOCK_MODE = "Continuous", 
    parameter NUM_DATA_LANE = 4,
    parameter PACK_TYPE = 4'b1111,
    parameter PIXEL_FIFO_DEPTH = 2048,  
    parameter ENABLE_VCX = 0,
	parameter FRAME_MODE = "GENERIC",    
    parameter ENABLE_SKEWCAL_INIT = 1,
    parameter ASYNC_STAGE = 2
)(
    input logic           reset_byte_HS_n,
    input logic           clk_byte_HS,
    input logic           reset_pixel_n,
    input logic           clk_pixel,
    input logic           reset_esc_n,
    input logic           clk_esc,
    output logic                       TxUlpsClk,
    output logic                       TxUlpsExitClk,
    input  logic                       TxUlpsActiveClkNot,
    output logic [NUM_DATA_LANE-1:0]   TxUlpsEsc,
    output logic [NUM_DATA_LANE-1:0]   TxUlpsExit,
    output logic [NUM_DATA_LANE-1:0]   TxRequestEsc,
    output logic [NUM_DATA_LANE-1:0]   TxSkewCalHS,
    input  logic [NUM_DATA_LANE-1:0]   TxStopStateD,
    input  logic                       TxStopStateC,
    input  logic [NUM_DATA_LANE-1:0]   TxUlpsActiveNot,
    input  logic [NUM_DATA_LANE-1:0]   TxReadyHS,
    output logic [NUM_DATA_LANE-1:0]   TxRequestHS,
    output logic                       TxRequestHSc,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS0,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS1,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS2,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS3,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS4,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS5,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS6,
    output logic [HS_DATA_WIDTH-1:0]   TxDataHS7,
    output logic [1:0]                 TxReqValidHS0,
    output logic [1:0]                 TxReqValidHS1,
    output logic [1:0]                 TxReqValidHS2,
    output logic [1:0]                 TxReqValidHS3,
    output logic [1:0]                 TxReqValidHS4,
    output logic [1:0]                 TxReqValidHS5,
    output logic [1:0]                 TxReqValidHS6,
    output logic [1:0]                 TxReqValidHS7,
    input  logic          axi_clk,
    input  logic          axi_reset_n,
    input  logic   [5:0]  axi_awaddr,
    input  logic          axi_awvalid,
    output logic          axi_awready,
    input  logic   [31:0] axi_wdata,
    input  logic          axi_wvalid,
    output logic          axi_wready,
    output logic          axi_bvalid,
    input  logic          axi_bready,
    input  logic   [5:0]  axi_araddr,
    input  logic          axi_arvalid,
    output logic          axi_arready,
    output logic   [31:0] axi_rdata,
    output logic          axi_rvalid,
    input                 axi_rready,
    input logic           hsync_vc0,
    input logic           hsync_vc1,
    input logic           hsync_vc2,
    input logic           hsync_vc3,
    input logic           vsync_vc0,
    input logic           vsync_vc1,
    input logic           vsync_vc2,
    input logic           vsync_vc3,
    input logic           hsync_vc4,
    input logic           hsync_vc5,
    input logic           hsync_vc6,
    input logic           hsync_vc7,
    input logic           hsync_vc8,
    input logic           hsync_vc9,
    input logic           hsync_vc10,
    input logic           hsync_vc11,
    input logic           hsync_vc12,
    input logic           hsync_vc13,
    input logic           hsync_vc14,
    input logic           hsync_vc15,
    input logic           vsync_vc4,
    input logic           vsync_vc5,
    input logic           vsync_vc6,
    input logic           vsync_vc7,
    input logic           vsync_vc8,
    input logic           vsync_vc9,
    input logic           vsync_vc10,
    input logic           vsync_vc11,
    input logic           vsync_vc12,
    input logic           vsync_vc13,
    input logic           vsync_vc14,
    input logic           vsync_vc15,
    input logic [5:0]     datatype,   
    input logic [63:0]    pixel_data,
    input logic           pixel_data_valid,
    input logic [15:0]    haddr,   
    input logic [15:0]    line_num,
    input logic [15:0]    frame_num,
    output logic          irq
);
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Jku7l8SDwt2MVSZLLZRgWaZSe46wNnHzAbbsBAmai+0sWryJsgSQrCGjRRLI/Bqj
xTgDh5NtSkCEjlv8nSlZWxCs53odOFp115a4d9S2JHJHhZQfISQXzWJZtHvy5cr5
LyseaeE/LUlcnPu5Cat16mkVY99KlZgyZDYF6kokbEhPsaHMXzEx2z0SANQJNkTP
2CW8pwfBZWVHd8R7+eghme6YqEzoZabFke8bvinrPef5hjI2vcJpfZZqryQmr4q6
7QR80ES9TZGp3LpboG8t5E99r9K4ySKS5uy1JlEAD9tBZEvqoBAO6FDYP3jWbwpi
ZbvUUKZSXuy/YK6SEgttuw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 21296 )
`pragma protect data_block
wqnMPSFcSw8xzJ8deahRq7ILFLWvNoteXW1ZxEfqjv0Url6c5qabppcgslqvrEVB
YUbJNd3Cx0eDp7ZmKtcekkGnoUSvX+XVL9yFEV64Rz+g+nLKfj3nAuik5NZDpsjC
DIT+ysXOqZxqTXIXaVkm00FUT6pQYUyQB+hurSnjxBmHxyJP0jraXL+HgAPcqGTi
/0L3SGbXFQ7X/qYugNdRo746lMtCc61Yaj935kkqGs5hNDc3obuNcZh2rC73mveL
T/FMoD6G+8mTitzj2AbuBB4F3amQVaBLbTWtHWyt7H/OC7Jl7Vp6CcdxdEcond1Q
PH8m4SoJXnpoHPeYJ5I5/QA/u7xa5ZgWf9gC80jAxEB/jr7khx9KGrlzFaE/iCY0
8iGjJHTQb8vvA5njprgP8oLUS4k5x9PNgIEUgBm/UsV23r0r8kbUmJI58zSCdYP4
HVXQf+VJmnb6xcaYA07AEEZnJy+dmmhaVZHFZ8IjjRMNmY0W09Z1HtNktM0ULVnF
nZys1Gk0f+VkOmqYkrJbKIsDln+qgpE+YosWQ9nqITHZBY3K7J5I0RFBprdatmUF
8T7Bx5G+myLW6Ko+6QuzwO23H4+YjTPXs/4+NbiR8MSeG2BxDdNIc/B00qG0ZX2U
RsJR+RSquTGO55gOU9XDOIvSoIzjwqqW41UAg+OMr4rblOduUu1slUE8sdnreg6e
k5HS3OHIJYzHRPlhXDTNOaEGThm4P+o7ylF7QdyHYdXwHxUgSbVYDsC+qVgiQbY7
WfD8KLyZLBKPag6RyDuMegIe0EEdUqI7ls6K0Vu6dRKjXGbMY2Gk31rBblyNsytN
V7EhNsYO4+DKnaAFL4tiG5T5baiKWvtZKihj8i6XVRpFRZ9N2Jh7XofjVmQYqx5d
9KelTWreKY0oSd8AdH2wXwpHqOgamtL0mexUeDd7fNzNeLgTSK5+2AnauNQEx5zp
0pNgESiRhoMzYlGZqq0nzPh/rmjE2AsMpRAT7OoobSVara2HYxN8xXPImOlCZcXa
LpZzf735ciC6AmKGHmcIF0tH+xDGXaAZgjWm2Ye8V4zQpH9jRHoPNSkWH6rBVKpy
tcIpUocg/pxjjR4bmvlYS3VZJRGb3DLU8f4tZ/trZurdmzodGDsBFdMxpl06tsNz
Gq4cqDBL/0bgZC9F1lF2H+fwL/MQuNbO2XKQxgJhs7YCbikRQYCSa3mts3BHCZs0
GxGxM5WRM17zIcNgxHLxxi44NJXAVc+gcpY3DQ20lJyFS4DanRJpS+4AKEFb9o3c
xhrWV6po5PX9XbAvZa9oEi6SutqlRhhV4IKVONAp+0VxVqXGReqkMPvo5eIItFdz
JeEe2bZd7mA6MGQorFZ0Acwmc/jFGssBjlRxaig9pjBHcgkwXxnhtGKzmvHk5XX0
6ZS/g6L69cKoK2bR7Y92YmlXZfdDvj9JlnIBF2b/OhRxh56Uh9TDVaWzBX9DfLVp
TIEVEJdd+zWU91xRfJkEl9Qct3k2ztcQVIPU5Ghq0yL4mS5u28O2bzfj4BIuhCF7
cb2kdU3b2+1rq94J7Ik0rgdYQaoq1YSKBJw7OGyXS33GMefjRpkGQTrIigHZnVjM
h9X09F13245Y314Ljos546kwXJz2ceiN8Yj7it5aKhBhjvFkP65tsRAgcr+atVfE
ZeQ+BqCiLoVIe1DT6MZ/02cKtD3xt6sAS+b6/DgQi37DHdhjrN2qgNtKqOrDuWvY
Gs20/NfEX/b8zP3hbfRzmNk3YwdbWwQs4nO//dwFRjZttOFEFWNCsf5u2bQ7Y1nu
bER7GDZ/LBU0cISUYu/c8Jbs4HUmwFZEHXypxswe3xprV9Nd0UNNcWJGWxsxWJUJ
mUTv6AF04Iv3FIXYRQpEaW3OUs13aGmSplcHH8oAf3KRXdmQX9sYgs7LauDxUch4
tWtRJJUf3KkKxloSaf8hpMdJGWBqIP/hEAwLzR3cIMz/mQUKO33c3jqkbdUfKgAH
OLzB/glH/sMdvdrhObnzvSaJDmdKeewKxR5mBtWmktguDxZzesDeMv+D0SRn6Wr5
pKC0rMhwj3CrDynHpQK/DZKj8wN+hS37CJIIO1Wa0RYH6/GcXlENK4CTosPZnWQK
pJGn5LRttflv5hbaWlTQo2rjTnX9v5aoil4iFpG0Wd6j04xxsB4j46vltEQhxrqb
YqFijb0Yr6c1xr/poD03C3SiYWOKwt6PBCDyM/kXNw/4k/xjjkpg5enaysMmBcWt
sX6I+wIGgzq1z5zbv5Nexzt9prumsnvFFHE+PBLSrqR0tSbg9EQRsPDSZpsRWKCk
ndWk5VaTFe3V+zkEOuNDhzPCSwwKjCjsXTXI4KvFhhZ1XlB/V1n4EDhFZn4VEBPQ
4+m6R9mq7Q8BsjOH3wyyE/c6aQMcHqxvM9PdGOOxNlxqo/gO/r3uRNZnngCTZv6X
kKVLGSpyy/BhYV5ipPQu6e7Ou1se2JAzfxU0VH9c71Yc/8VStdCX04M1rYvxixXY
LaJAWZO+e8CYwe+oC2vwLRHx7doMKlWW3i8jNv7Y64R+rtaU1JcO9/wNr/xPAroM
uRhnsYUz7yEb2bkDB/jtG6lwA2Q+FaTnJL1aRZCsFFQ8qcDHCG0vbZ4xla7dcTp1
hAPU3CFYDDnp9gITQMIRkn511j1b55/tyVm22LRiHAB8QvxAwi+yJMs7rlHipxv/
1LKMu3JMpDF1G/XRvwO4rxeOgInWm4th2IxuS4UzGpbFQZibKirP73zx5bzO3F1Q
aBcCJbNApUEh7WU9pTbvT3QqeKuLsDPqlLcFkW1DOWzrr8ezpOkbNT7eqq8c/LN4
L6ycPzWGQw8zurmUDmXylNO8DP2qL/WH/LPOpZvVDniTtILpK+5zGZ7n0U/PYBfO
Fk8L7UEwl4E5YhgL0TmrYMKMsfvw8MTsGHWK89ZEkxmMoPs6t9F6h3eUU47S0UlR
sIkYrVmTezEfhIPfNAxUu6Ifej+o8W4z2iin7V8r0xhElYnZ1R1GusVTO0kZgUbX
1/gY+YYroKSXiTbP/Ki+Ho3pL9btRzpkLfSIgxtXCjWK5Ksi7TpYdyxhD7f6j/If
0whMm7JnNTFRbSBGU2dtqwU/HCxemB3Z2dPBF8eWmYZdvPFCLdlBNKs8uGwHXMPh
f7vAkVSq4rQzfKdExkFmMld2RFrfxL+6QRzhn9rbWHnAdcZEOMFaJAVLEi376qLE
o2Wz8XAOIDP2tHwdVepwKmMfft4zqlbOUDPoUHo++fSEcy8Bl2GzA3OlJTFaXAb/
5c17+Y+IFEeZ9GcOb0ToK/HhaGby5HrP+TxMjwfhCuFPUM1Wxz+fDcD1ighxYzl5
qNaksJmJXDf5bpX5zZG5VaVpp55dF/8fbp9fiij9ZhOySlfKTQK6i0W1Ej652XI8
MXxJWALktbcafNOEixRUYYwUeims1WrLf6RklfWeZYEbyxOnxMNJzyHcwd9nh5zN
2giNWcY8vGjYjHk7qf+FzsE0ttLjoyUcbxvMx50uJUkxBQM8ZF7BZr9cbSJnN6uU
U/jormAgbCKfkNOykwiHT0WX/jIo2wg1K70HTXQ11cjZUznZgDfL5cP77sCP7mtE
dIHiSC3F3iFvfBQTWACT2hX9iCV86Wi7v/acfOK6MsuHO/+tjQGb6hCeur0pa8uJ
80NvmMLkvg7JT9cQQmNpk+9Ht5oZ+O0SuQvr0mhE3BDSWygx6uenwV9Ycwkg6DtJ
RyVSpdLHVhrq6jSqS0sIVAPkScqvXbswi84NgBTUiaVXqGaHtL8iABrLNsc2bTDO
t+LDQZmGjdbtcDltepWaRJ3eFOaEVO7SJjXK2O7K+caXfsk1O0CwpeN3UzSzTCcF
/wz86rSRmwCe5AjkZyBKT48Gb93dtENvPD0cFuguO5RVBfXFMeduUwgqVfpegYTZ
ffM0dLc+C1YmNyBrR1q4LdxGec22KzSo8n0T+u15w09Mc84RjwVJnIuLG1U2NnbM
9FkScAzcGdTmu3VOud/oFdestPXVyRBu2GJtgDcnIdLgEAE5FX4KmaeFeL5i8kLp
PjbZTeHHUG+ed5uvnFWnOVnCvmOJ3XZcdvT8ip2CgD0kZRTVo9Dthng7BVwQV873
8i+BkYrbD3zYxVFyyNDW3zoxg/5P9f+oYQzLu3hNA0P+g2p4BtU+0AkGjfrt7MJ6
C7bCb2GQ1lSD4MxaFpM0aARcMmWY4Dq0fL94d7sSYM5OO+nBp89UOrMQjs6bGQ52
9qsob+kfQX2zhxqM1tIZhxw6LLM5VGmMWeIBrylbjGXPigK2W6LiQIa1UHF1XYII
Sw9+2tk/phdBPq2kyCFlVqwGmhcFlAvrOjDrsWotFap8CaMrgWD7CeHVLfDy0b9e
WaX/g4Z7hQA+AAcPPZMuHyLAf+3JlHDh+hjdry/OY42UJ/MDBxuHZG1KCxaRQOrZ
61kLYJo1/rNrvwUdyNZgdDA3j1rqTYstUZ3S3DC7Wggc798PP3VuO9cW6S/Tzrr7
bU8LRjGjH2lAuR0D9kcI8CcLqsgpBlk/+d7ISbU4rT/j1VZoHOvFvVrK9gPNBIVR
EgQrAl9+LAanI125onXGNtbtBxl9pCc5GKNmMnCnIRPJ59srIMLS8mG02+Eigcbj
PgO/tXaVj2FUDVT9Ox2mp4BgSBjcwgNHQLO42iaoZqMwWMGJZIe70/CUY+75XI31
g9aIAr8spIQ7UDTFY5VzYDJc4OWee6vMv//Yz4RJsM8wx6gNebXuHUcPIlE6auOV
qfVv0edcRHe0UyPtTum37KAQBn3kQlmT/ZZr4Pf4spcNkUaN0EdAwQk6k2EysJmI
NjXpKcgcmmGhTS14E05wU2jXmdmmJcfkHw2BMzTOWEmgFqUJkd2Pnr4BfDAyXHhS
+0iwn3Kv+yC9m5o+6QPMIEXB7rRuhbbL13qVP4TcWuOHX9HpH2LNHw7uRDJsIj95
pt9J/w20tboyw0j/yD21PCRf2N/jhX3+V/5lGedcFyEFufVLehQIvTRgc7GQu5Tb
cBEu+gRwYeADcCPG+T+MQQ0AY4a9nBrFhzoP8So1CmCm1h5URzc2d0/JVclhANa7
dhWfLGu5DVeH5R+Vai8JAgBXILYnj0vwTRsE6JowWXwNAuyEtyKhnwW3MQeu2BUX
QAIknZg1dNUmoVSOefWRWWQtPnejdzLnuRsL46U1VLB/l22W+UF7hOjAxs8+eUOF
qySPpuwzakOgsOV5Er61vycBPQyZcX2zzGQScM7PaWNlsQCho5kNKd+JgfpPaDwf
oAj7woNrjCV3R8MsyYAPY5anVZt04x5enBUtdBbtAzzEaOTMP8XDAcKeN4BLnUob
yAs1zFruQYHhZpSVYjbU/z1aWEmxYB6p+rMhDSJj2gyhyPtTzmD/lol95tttMakG
0kbk01t27iaQUSBsh0jYc5rridomvYyHmvzOs8kOYDD3hQB0icSP7aAEpZ6djAJL
ROPmuN+Zc+Db1DO2bIbBwuEpsBFopzd8aDhMFC/52tQmoAMpwao3rRLVpvL/2ax4
wMywFxBiZPfQTbb0OmdBn56PxQ9rYsmD8vi+cYQOLwejdiQ8GrQAEugYw7+cDEZx
l6XiiLWKVlmegKQa651rvRmN6ndOvnwzi0d9Ttgn6DD8+uQrmqHxZSc9pWmib546
Xmt/axJ9nNhMAARF5NAe81fHvIlxU7hUksvDBCbREnO4/2G6osRm7xg8YONNeBZR
VR7DfcwI722ppgb3dew7IQ2fzkWAOdeB4SxOuRNGfrmCUAqOzcuOt4N9pJBLDEeI
oO/kxgCxV4XtwumGeG4hRO3rExNMm/vGbXEUCgYu5O2o3U/XVnWASsmsc6KNJnPR
1TYtw1noPomnG7EoN8YjbXXn0Ozjp58fgCEzYa+GM3gSm0w2sChVpBX33MBng1tG
WG6Mgii9FpalmZo5s6Lt7/84IappNggnBnCQ0/5GhFH1XC3GedSiPcGEyqm2xEVR
n2hUkcTdmAbx7QZjeQ5iEyOG/h+Ek/9R4EcEKcbMJTVBnqFuMrr5fkvC0rYLnA6H
rWO/oTYTgtuKv78QBn5LJEi9L1pceVmbdbQ3DXhQlRAE5TjeahmtUpkfs1sDjABz
1rvnxX5iw4Dl6YroY7W0ARDhf6nIbgOI7P+80W1hllJZ784Vj7eCQOAWce+7Cx4D
XB4oL10iuzQs7afJw/f/8pwQv1QAvjbwSuVZHCbgv3yfmBQI31orgzgW7rrxAPxG
8fMn3tA8QYhFNSMtN/M2POKwg4HVb/VfeKapmt9G4JDr59/Fu83OI5M6wjP7mCoF
MpOas/pjCjOk0dC1qNI3r51IK/YTb5fPVp2IMVAs77BPsKEGCwHSpxuEYO7RUiAE
uvEapRyGBx4N61851d9bF4jxC/k/zHuMDWLC+18o3tP8/mbSOwOuULqR7aR+3hY6
PuHEmdmwrCogbf8zmYX0DqLVtk4EyUvY4mAhcEuV3RLoEyxaCUL6mCf2fflxh1XN
vopGUp0OL4UGq6WlXxmZO8E00+L7MXWj9oCJCfAVCw8FxM5Y1uo6bJbkdYzxkP1k
XQfF+ADjes0OpjUhWZ4jQLXZWzOW18/+7l4IDx+DbxaO8sk2M5lGcQQqLNTu0WKX
x/CUYSLKG5JDKJaDBpPA+9EPcPX7G0Ci2AgsrLpY8SWWHctmXxUALGXbqjFZSb0m
rbSVUKJovAAlKEkdyZg6gCMMggPQCbsC+kygwh2/rYQwgvv0yibmrEQDwyJOFSHc
sfWMIMo5Spa8wzfGgapCxMVO9Pr4gpQJqWVphEsnWHyYhak2B5UO7vngz4aqrUyA
70I9wtNyOut8NKSwFYyfvl6vNVcV77u/P3hPc9r9KKQhhe72MVWTVr6BtaSa22+t
plTaBmJLTrq7JEl+fGrhyKIjVswh0tqtKqPOGbzA5PXQ9ZDx4Y2JPRj4WfTsMK7K
7lcq3qBvnMOhS/qTi9x8RotNNMxwUaHWC3V1qj0VWqNl2Sf1kLD9JgbxieFGItv1
m6/7jTHENv08EBpAzt0OeWtglFUZL+MbYyLDZveCIs0WoXHZXGX+ZLAapV76Cgv1
+TfyZrR1Ee/hcBjsZjKpMrJ/a+LR/1axqpk2G3qM5fiLV029Zgz+m2ZCMClponxm
VuNfdaKv3OcZTLaSBhmcf/2xvRXZkY0c4FqPnnGQrr5+vUvc8EExyBGvIUPUtfwx
qSwpgQ1+3sn6o7sWKkKNToWZPANLb8+F/j3pKgpiePw6/o/h2UE+2D/ymldTsAYL
YZifb3zhOU4Db/Ojd7ge993luV9aq/wc3pGV6N6ioGbX+dny0mxFLcZ+3zhgR4Ri
R9ufS/3olw5hxYJ+oVwdnwnTrTKUOsitxHUFE4KQC8vBAfmGinBSu6216quKMr4a
6I7uTG72yEOz7pz7n+J8N5/jrScNwudFoeHQi7MKt9v7glqSmSDPRaZ/weCk8r5k
5EfvLUohYtV+cjFRGjnTNnH81nLbcX/9qlVGhMTDc97AnV2CBP1ynP9x4fydRuJt
Jrsahj1U+izSR7H+yTuET/pCW3PYDlQoo7twtIPvL07uqqHqLtu5jBJowPDDrp3B
ZlRvb+zj6Sp6530ja2QNTNF5YNu9VNSsD3OiwoVlSfjpAFJPpOArEtXQ8r3KKx7c
NQ8yZ0AczzK96cRBm6j/3PSo4jwUFv+zh8wTxQd7ReB4XN88la5FZUhF4ikfOwwT
s0hXMoYoDbueykHCj+injHs0tSbC2FFIzWPjS5OfozmKOvaKM/rbKJQJ33XBRonS
SbVG8LZ/2CxnP3/GhSSwCCRlccdylXd1TMzQJOaPnw5l7g0wLZzUWkbHyXiLsRad
F63KILe4G0fym/oT4n0nJGJOlHnvw/jyypIH0SgzJkWd+2mD+hIhWs3bw6zKZTRG
iHCE0NmSCt5QcnpIfdHnpnd5cMs/NclYqaE7ICNrAh5wXmD9VF5qDjhMy2IpqXTc
T5TE7nDGo6CuFLpBnyA3HSRzlukHKGp3n65W/7ZOpijzLHcPal1xQKDMDyypxOV0
dlEPUymFSkfuAuET8I6Fc3+DH8/Iygah3DG7f+XzjcY+o2yGK/h0G9EcuHmxD4Yf
oRuAFqt+0tUCmTLElakjfonfrWFYtzwmDlUuuGiA2qr7GPx3BnEMROUjNeHZpio4
W5OwEY3YDHDJurbtWBg3RBjPSfFUwFVU+N21xmKUCNUuXW4WmZ2EThQF1ooaQkuZ
iLRDwOiuh4xCZcqNHIBcwYzFzuW8C0CX1ZOFUNKxEKXcfKUQ573mfi2NzQMDy6mH
mJmfGJa55JL6hl1U3RD03lwNWmgofvX8j/umE0nDRs9fD5oxiuPpFN+eVvZVF0xE
fuiNWdO0T0QLJ2TjDVr7OYLOHkwVJAGR5PMY3MGBhLi3Mb2fbtOM7DSZ55hIE6IC
y916Ocdg29CUh2RpdImDMnXE3qLW58b1sgy3D/xP76PPWp6PeeEVO+R3skJ84PgN
JjCniQF1XIbUsPD5ugG/3hQMDUMujvpI1wr/BlAcHWTWYYiW4vO7SLcUscQYuTva
/UxhEWjbc4CerC1PuL58BGW7QzoxsinW9eDzXA3x8Ok6UzVzk2qbtVeKCs3zYEkc
+3K9OyhohfshV0/vNFr8r0/nvc11F8nLP73EtntXt1BKkIs+odju4MHyjHL+9zlq
Y1xFVQAqy+fq+ssE81KjLmM0ndJfYru/8uEEETmLguDlT/h5QKdhD1490tdgAQ6k
ZWjLmnLxwBpsoyP8NK5f1HRma+J9VrOMXu0Am61nxeBqO62AWxQU5xD3ZqQSqNWl
ingBQksQZeGW5e+XyR51kc+2hu46HX9J6N6EEdG3YCQwOAfZlE+2QosRZJkNaA9Y
05H0jSPimT4TyYt9EZRGNmU+W1XtgtiHlvmzsLxYWOPf8VVoDpOSbbFF4bWltNQX
riRWudxORk9oSFm1Fy4m4HXf3s/EHqUE9kv6yPTs0KrtZ7vzrm3DPM1QYeCjK2lj
SQ+Pq/juJWahYDp60u2KS/5ouXgqIgVn4R9cg3OnWwyMm7Ljzsdj6UWJhTpTgubW
tTHr87Gvw6WcNzjSFs4/JEVkmeYfRlSrV34pK9CAwbKG/LszG2A89A9fo7/4ZcAx
VCL51VjX7kul5CE7coQfmCSydNX9MdPEyB/eJn9kzuqWIy6WaDIZ3Lmf5WMX/sBT
czvN551C1pO8oOHQpbBrW5Rlrw00IMoaNazGQEY1AQpCPIfqvJ7VAuMu0RkotalW
lrYth5KUMuQoND5O7cM2/D2KEi+9G0hmb+BvJd00jN1pmD2g30UW7ixZqTsAMGCV
ED7UMtKvp+PLHXaBN99QsaS6KgkATGfc5+WkZfSlK/15SYcv0Mq7GLf/vv3myGpS
mv6oi7c9Kyc7QyBoyUPeadD+pJUd2yn8W0hfGZd5aTxoMVMM9iH1SlS12nbBoP/X
XTMgGw2npOim8kgspyc7HuMOKZ5dTtHITKOEgstA0eOH/vh8yR31uh95HcxaJy5c
xix3Z59A89eARlD8KHR6KHAILJK6u8Rw6kml/OACSzNuABTY91xi5HgMxuY/ihwA
fop9htvcNCxEUWN/gYaBumg2it5hg2Z1WQLRhvGX+nLFlrjmibNbD6am8x8Hil9J
7Bd2/4kaIFQt+Z1y/RJtQgA7ML8XbiK6oiL64/IzJNndNkfrgDJA5u/xxxwirage
iaacgs0kyH1ztKSoVDH8rH3DrG2dohrS3SZKd+6qLasIEDZxZwQjUH8pOiL86jm6
0FTeaS9rV9YzYG1JEF5Q/AWx1SJnIeeN+rkwmGHvFHVSl1LudnpkJHsSaA4CN0mJ
myAzfYOsscYuGX6Uas/rZOHCUJHmcZwiymnFcJI7+TXq/EeMefXZWvdrDkJo5/Mu
uAs2GBhwJ+Q8Je7hh1opnNkWkDcILn8EwH4ag7JD7Fg3HYZoddX+rxt3MzEyPneO
I8k+1uSKJar3BWuxKL/7ASRaW/2nCNQIfTlEo4ZR5AmEaxFw93m1AF3iNGpuf90/
Ly/PKp6aTakGSXJMsUwgpam6WcS9l77mwcnPQQbs5jpzT1pygu9O7zzyQaK5e2te
D8mR+qZugLMTT/VFEXD+f3Thr+zk6pXtHKh9Bjfsq+1iY46Rz0PvfjHXsuvtyefV
zUGSotekn6yhFjeFC1iGapcMisg7NE6KfNQi//ZpbDbviDB6BA5pvPC3+OptyS0b
+kDONLomTuYo6rDir00zXe69tHTIbLaI6XIrF7ajqgZHdMo+p5GbniwqIBnJdysl
muDC5nH9ZBZOs4JfSKFweTs15no8WSCIASq/Ph6N/D8mlPQxUjNv1ZTogRVyyQoI
h4kRQ4v0SVe4O8FcAKd4Ar5zpO5cQhuwveXOH8+fgGkRLwtPWLLMXfQW0UGd2SlF
Ds5hOvAavv4O1RUT3fHMJyy1Rc1QqY7+QTcwVN0A3YAABy/g5Ct5zb5pFY5cnySW
Op7XgPKiP12s+jii6wB0xrKgGhww+iS5dId87Gsqg8kpecAJGN1maAjbZ2dGx1wR
AGsQTmZanqJ4dzNDkRG6XqUB6LvPRaCOCe+jqJZHTqWZjSLaQInCXyTq+HLIHgQL
ZtTZTijS3wd49iSRUnExT4j8UWBqfdfD+vWS4DbeZqOTpkg+x0ktjt+QWU5+TM6I
G0GDeV38BB6BA7mR/pVsJtWXPpkdhmp2njwowT6ICjVV6eLUBqBVq7M4FKVa0QPR
NX/FK4PH9rV4jaLuGpHsHnAEdWOS0T5IUklalXl6gAzLNIJZkNV23DRfzNk/1hV5
DC7ojyx8rOW8HyCofwe5196VXJVp1sLm1i5pGf/1nW4aYTmEte7nTLShW84D47p/
TvvhWTVPFJvvN1TJxsGmZ+E6cx8DwsBnRRq54KXkFXBG+svgzNR6OFFDLS1E+pfs
pHErpUKGXRolcZaPebXNKhjtwJHe4Vy7iQA+cqfRSqARkcWtsHx/boXB17zNQybS
wH+cF6+tetIwmldIILnpy9MhshD/P2g++NIi1rhNvNzCT7sKSxMLLv3kmgw8U7iU
M8XOtrXtOq4FOBP6fZJe781wX3bX1kMXV71H0vXAZqYCPp3LP4zjW2E+ZM1DJQL3
tq7UqYZ6ZtkGF7s0rk1N5TTYUjZtt0YPv0WsCeYOojRcawE0YkNVPylpLIeTdSL7
H2N5UvJQnT5e5W+jSd1H8kuP13BuoPt/8vrsQ67hfmQY+vaoMWkiLuLfHXMNlFSO
h3uaP5OML5m1te40HGrBxLL4pS37kxchj/XaLQr2Q4CDTQrGd9pCfAtZrqCkvwP3
pyJbd9XhyOqq3+9X3cwnTWjBylKl31Qwz0iW1uBYNqBrXqXwE1wDQLB8Ax08lfyu
aFpxDgVS2hBij+P86hqbuSt3Ty8xPZ/siJ74JMqBXVzQBUOKEOWZdMriFKuM8bFh
ZX3en0QuMeprnP1DKqsRilNrqoNp/vMVmWSU/Em8YHs6gmPSlHeVXojCXWIREGme
fWckCrYbyKE4yo2fB4zfMCaEY4rcVwsiqDy/0ldGEhK1mfo1bIl+YoA3fUPvIbyY
PBEJ0kXgz1hNZ0b8suNc6ydKjdL2osuqXlc/gG4mW4578BerRRThZucjgkfyPgFT
GWb46wL797QEb85fftcQyxOL8+roFXTcaiBcRYOOhyIhKF1GE4HCP3EX4+uUZf8w
3OemaKFd5SC6XrvesJfa5d6+R15jFmF9UXTQJEQdxebkwuJIJS/v73+KurQNthLy
gPs2nJyhPXXlL4H62QKCb6/EEabqVk3HOzQKENCab9Pu4Z8rgNkSFYn0k0awWK1k
/eHMvcJAtukhg48xspqV/SsH4N5OEqnrBPdBfnqJKhtb4taN+KqKepPhBQpOptXW
8o+OMY7S4wXc7RBeHbxOeKku0SL0p/aCwr1LVAKZkrWMoW37JhW5rCgTiAnWRoO2
r7+FsI7Evl0IhxpVhHtHBQ7Eai6fdCI+Nfw2NgR/yZL9PNLRA2vVA2hpSj+dBUDW
XZQRh01LlFEN8HTjfXNPgRtZ8iqVYk0/juTqjERwWVYniTVKHFCXuR+4aPNj+Ifz
EFhVH0t6UFfCEsXVcmM8BIzocA59Lq7QlOAVIb2JjhsoPDX+ZJKh5YlRoTbDX3dC
cHEU2SKSEdvpmvSACHd+r/ZtltfmaKJdZLsBGnM2rFFIxRAQs1VKKteIeLivT0FG
Pf+brrY3en+ok50+bKqo8lVrqyoKf+YgrGWVHpCn1kZ5Hpng7dmoIxYdGP8fE/Jq
4Im9aiaIvrEpkWQ6kH6XexcLfngVnhN9xdWujjo3LRFc6x4+3zHqCZGxGgGyIBZ0
4Cz9f5JDnvldm2Qv0Rqf14nHXdB7yf0PZnerM0X8Cf1bO36NmD7NhuwmuMu4ZZyo
9s8Ayh3PZTiDGmKfSMz2JPva+9pA6HGLG1Y9yO2COFIg+HQJbwfNXiPleQDuB61V
OBm5az9fnVxGaQolxqpMyH00QedYL3X0IVj0UZbiRsoACGgKHIEftXS+SaTqH5nH
SFoBnzQb47ss8IT+8TlCCmD6p85WiqFHEVGQJRfZze9YwUF/EJFRReJss2V8l+4N
lQQq8rrkogTBFcd6wQPWcRzOOY5ixZqnMe+VIHjZ/iYur0Zk4eVnbsSXrtjd82sA
x10M4Hm6JXD2Gop9CLz3HzclPYEmwlRzpW+zdVNYEiyWQnY88N7+DIV1QahcKwsI
p/uTTGg/wOEXVheitmHToFrAfUabxdpKq/6UwZzVjD4Al3Zj6AtHoIq7jjrsHKff
KOQK8elu0g+imyJdW8bRJ0YR4MH1b0GramKGCHWzf/zBtgX9oilO4kjAc78Dezq2
IS1mIDsZRyKi8CH8iQ77vfdCCXN5gyGEsFTYIyy6jaPcLW509Xct6EkPPtwBxJX1
QZ9sOB+2Rmey0WUau5yA7rQiSHlnfx53LwUIFv0ROjgF+6geuIVJ9NUj7i3Yl+aQ
8blE4G1T06TJNfmbo9Z/kMtSGisLUrnsHTv70y9J/3mcqPMrYVuUHiFSBiKiJyST
W6dVc4yXLEZ+C+trhUhzM4EQ9sMAA7JK3BJozAROqESK3KHZ7e41MUmimGNU3Y31
JoWxy3wERxGioalzftjRUnPHDmgu1EJWUKrAC0vGFtvyevddwaJL4Dq490KnPXYJ
/A9Q8IRDKuveElzqZU5vJHPj5fdBlZLz4DOcJDkpmbVMtp6OeE2nH1xeo0acX5kc
mKlNNSWh4IhjpI3anuhmeREOZkw4BRnL6IkGi3fOKL4J5trwWPn+DTiim8cuoYIn
d7HpIGanSGD34Tt8OGz//RQ15nB+wa5szf4rVtccjvR3/4Dbh9V7S+KiconHUA5K
iPvHHo67mUhcQXeHeZ5xMlp3Co1tCmSZdzjmmiA2Cf2GFIInHePjn87Y18LnSDxN
cYWoKdcCdQrPCgA/NZKar3SCZ6eD/V5uRtvqueVh3j0xovdvoYcMkZ+H5swj1nh/
Vr2nPQ34q07ZZyjuV5ZX+CR22KweDHe6X9aoEOaxR0kYwL9ggxTICDN1iWD7/y5z
Xspo3osdYxL3TY4TsV2vJtOKOaXGByU7z6BoZlBF8m1TVYFsFKqAyBNFrdt8VLYa
ps6uHZ6MY2BIQB/5FhLWqIjV7Wz9C/WHDJX3OevMxI7dCKwzmco0tOeGGVFvaIN4
nleTBceBfFWMo4JgGSQOaxd3QpHGIX2KdVKkvjbQ/VmRtgz4LKsyJl6Yq/QKkhjg
KIZtcsweAli8oPAkAvkt7dV6Hlbt+OG60F5or1oaJqZFVoY37GiWqljOFSNDN9r/
n4juFIK55fx/LCePBy29+SyU2wxYTnnuOjVvyC/dBKm8VIDcOrHOGGbapkbCRjBV
dLWyuhyjh9IfCnTfNa04RWzDt371PG4RaahVd09ub5dk6DdqUY0w+Rsv8+wAVXbp
nWT0WB2g5BjaX58koYHdsbmeBmWqRqIYm+WcH1zJ5GXpCPHjPu5wS/VMk8eciHfy
G0cUMJlReKiBZjY9mtXzqmtXttHEjT3vxRzwW99Jlebmb13U68hfCwNDqL/x2vad
Csb0L562jeDt/EzTFM8twRClFWcOFx/Np8uaDsMuAZj88xHCKktmDjbVkZnvH4ZA
wyqRRogq7o3wvmyo8NI/R4Djn+9WOE/S/KfuQl0q/R/6hhL4VSBun3b+YAIlXIE7
OZPRtpcuMM3aW+wo1LU5nrPsgwmk06rnraWO9PByGuffXbiGqjyo1ZAdo3Zd0orc
/uywsLigjpaUoC3jrpJTj0wHN9Ueq8IJ3O/k4TJ82rd3hMMGoLmH75fG3+xjNT6I
zwL3EHVdQx7Ez7PuD2SGKFd7tBWJpb85VLexbpY8+7axxG9qgXFJCeXQbf3loVSo
AHNyHluTFYHoOapYNgFOoja2K4L9I3IBvU4Srvk6qPKdtW4jt1mRdZxadmT0eZZg
85KmnMMMT19QmTIFx90hu2DENJhO0kysu+9rBIVebg4oP/sZFzMVhD2L2KKpe0O9
4+JoUe4a5l8d2Xc3dp/jh9ZrggT+Mf+QHnS1ipCkwnn9EYp+PBoCnV7uyCU58zpP
6Do7Q+kN+4Bv3dE6q8IiXPaJlHcZHJh7tSUJ287xrKbjA3iWyCurGZZJ4iicF6Rq
R36ccYt3U2HTtNxVqiFW7unzx83AiHfR8jFAWRlSMvlkdjpjWn+WzHsYmZMESz4d
oWyFTAhW9sFvxVBlOeRU67Mgjq8GAO9HWF/Vy1Z7M7aEVuQz2RAPznIWG/niH3Nb
si13UBEPEtsvngaXpJZlN5Pk5r1uROAe9f1NMVCUVwJJLDM4k6aaC3xUonV7nF2S
vK/gYwEk8eivwzlzGNC/TQiHbo05jzaXzXj1GN7RWWFQj4AvLDOiMREb1ug3VCIs
p+vxCcev6/bxXQOx9NorTnsVdW/vfACi/hfTXaXkDzrVI+Feg8Wd+RBZa42XUHRK
Qf7No07HHAlJF0hwATlr2ovlX0ZlfgvY4pVkfB1a4P6z9p+PVPne8Ri65xvAAY51
ZP/2nBTy2zpc4J7AgsasBzTmOBU/2GqSGhZXiuXO1mON0JGGdx4tkE6We/dT3sgc
hGr1qgmzLKhHnheO5m7GYsn+iIdlTw+aMa/YiewI9W4xO1yqldLDaHcTWPLt561p
wy2jQdcbZ89WTsJxc8a7nr5/v4DLgrs1LZQBWZCn0k/oU77+Sp7z7IBIMA4M4tgj
SpdSi/9PkqnbjrzhDtbXHpqLhNv3z7zfzY+yWx/ZHPn6PZDi7HXOL81JihW2IVwp
J3JxTSZ/Z+QYVCOkS8iFObevSmY195+fai0LiiqJa0cM69hN2//xALAvIDoOLYq2
N6HnvpHZlFgRMvCWELf32v0S3vMxSwcuNJon2/L5KWll5XILM5E+r7KFYbQwHVcy
5l9ZfKe8aQjZx7xT43Y2AFrxy+FciM30qhWTJpM9gxW0mGl5pb7wd1L2ia9HkBBx
n0LBDWJrE8QjNAbBjBS7BXwpuX1XUy6QeyX3klpSZWCt/TnMMkkWgleyN3zZwOno
rdR9U86ozOA9+CndokgR8/vNw2pGGathVv2FbifSX0vHSVysWnIUUcRbV4s1bRY8
3ynqEaxKkuWFHO3aOhhgrcFAsMWjiySSPg0Z9pe4cpkrtHNAOMQ2q7a8bhMHO+pH
Vjpsp5JywaZCaa2DruKsR482jZAUw2eFjLgLpOnrqZ01+E0pLNldYeEzotpnQX1o
c2Dzq14elLkZI0E5kDIUtzgrFhdVLwHHCkHACLECnnsRR3GC/HABQT+MBxxE8Ak8
vyBPJq9LqqmH5f5hDir5an4ArgzGGxKdmQm0nBbaaPTThGXQX15D8uzuVBd9W6Mj
FZs5Crwr3a/ISWK79pKJPeqH3JXNpOgNROXzvj32oLbYEHCIr7PrY5a77ceSvEeL
cxJs0M7u99O9QRBacu8ik/1AeJZyB/z4Muwl1rG5kgr05fAKb38eFS7wAWbEKDtJ
x2XQ09W7t/HBcJAcniG5qu7Y9d+jV3ze3L6wHW+WcH12ouJ2OJwHuYgeF58KEmPd
UN1LVfvAupySd1suHexcfBb5TbVCSl2kBkOJ2q2VHlEVbwVG78bCeN2PKOzTpozR
orRO+nyh4EJj44nAkUq+v2YDH5MGEipDBbApfbOq99dqiJfr1LeYNqMX8D5F19v8
yKzDBI8UPN1nJJjbqsgYPK3vdNuot7iA93fBmCwWpMvYOoRFgsZfwhdJgYbX8w9j
xig4TrC3uiay0hWHWkaN7XvE7guzItuIul0qd7YC2uZYfc68xwf5vg3tYyB5ePSC
n0ocw3ecKVDGgfoM54PDJDCQPi5gWyBYZEtUwkK2lPXamkeNiXxUsXPoJUM6YBGM
VY5CLxQw4XgbzQjrieE0CP5R7ajiS5xYDFL0iXdEUmtZyF02EpgT0/3SrUxd3WKJ
6Umb+Aw0jsgefEottfDNaualOKQAOzVDFCYoZMoJm+O6e6ZTcBH0Poylc2osCQv1
Lh04ciDYQFdBoTeqb0HBJlM53WWYWKzNc8Yagj0s/ufvw2FIIDinHGYb63hUFiV5
Tz1/7GDKDafTu1nfXOfszUEBAg4iiY2zla1Rosn9hxQL+J/yl472FjeY63xzB+/4
6+HOGbHm/ojB5j/DGGkIh5IFUi5akbhU/wNc3x+jsKvgIR7JPdRjs16no42G9THt
f/iPfby+QQRPk4qhu38llhCH/B48I5PpqmYR7+kC9qckt3VG08nAYxqhrnYKbIRQ
aE+Qesj0HkRLJSw5YJ9GBcx94B3VGFUnbemEOLnngp35DW7KhnmiCvEOjw4rZCo/
c/p4gi0Cwy7KKsUVEANUC0BHRI0aOGfWEI616+W1MLrq/2UyqNhfn80NJftECPmK
GCoHZmRn7T7Nm+Cq29e1S8fGiEBQPjsW0I4XnKbmkiAB/Vc0P2LvFXP8mH3Akb5S
KH81FAAIMzwW0R0WBrKk/IMqab4MQOj6kQumHueHnEdXcXcfcLo6VNTEcFjnDDVg
zTtk7NBKJThSiBg018+79n9Syla+ARZqrVTplmxrLlodDyAyo+cBKKhMgKFUNdb4
S8FQpy0nSoolaqHBhIq6VlF0qoUpRzvYbZ/vwtlbhSF2+qIMtjYdRkRsnFbGD4sq
p035wc2DNQS/3+fooGXYGJBLgIXdrUuAB/25w1RqhPowwB+zy9gn6qtyt6MYxTe3
sKVWxmxpymcg7tWc0dTwDcYk4M3XCh0F16ldGv1A6kIuRPH9jZWRCLmRE0ejgIAY
wb+Cai5BweapcP43/3H+at+PBOOXgNyOYbyHy0pbF2m14KK2ODp+SDtz9qpk8XlZ
62/7lCd08qWrZpMrHIk9rGGwAUBNPgea3ctJtD611Q1CA4HhhcaMfOlWTYo1uipC
CPyTphHSD7mw8M/eucmojMP4kad7unYXHvEaXvT2H8cFgTPB/UbLlERBonbwUANj
qdnsuxPjCDWf7asdL089mVB0O/y3KJ5ztp35rdi2EzodtxdaFHnWbpdgmwz94yKH
m/WI57pfuDMp7zGe0cXKROZFlb58NgxKZ/W2iBuMGALu9qVnwMv28TRq2aIG6Df6
7y092l8TvRojGuhrSLPKBJoNtih6Atqwu9RmWmcTvs2dqULdAgpgk4UovLMySa6K
FaWcItQuIadaQVpaS+8MFtSwJiw/gqMEcgnykdYunDsVe9bErKbcIDZJ0JtVL9M5
syj97IgoIa6ZhMZTLSrgm+g8K9HObIxnx2jECZ64B1BTFsTdDIKYG409W3Tgtici
Bn1nLCfcPKgkOzreE7H2yl7zYimrpkdsMJX4J7OufG4Loaab8MP21sZyOURRhunX
6WtRVGqy4oNqhHMkfE5JuEm7pBMhiLR7hjMvt33j849YcKUA7wNSLtVppPT1oMjC
2Mj9rfOSYBxk8gWQp1BrOrI4d/z+rZFTWkYFQ7Ip6ZDbI2e90ztjH1Jfgt6LSjhB
fdKvULKJMILRaJr0zoX+x6Uk7bXk650Mu+dgvKIHIXUcbI77t31oNM4yOEOYtrnO
Jze1jUdpKidYlyptwJyalmLs1+OuCOYqMxhPmITbKW/ozb8HiPmelozxJ6r00gg/
oF1THHeXlmTAyrLSJFeHTHp5Cg4709tGDhgnjGmDrXbDJBRNxOkIVo8y8P0cR31/
fAGoN94lAOku6gG+OE8CuOcfsR/YSEUCndf9BCaW8+/WlmhlmvvpfYKQl72GHeaN
uCPZlA3H4Ov8f0cfAsai6G3l5kBKolrhUgYysS2SUzbdFAlHUEMoXO6CuU/aMsbE
WfJSKD9/x8WdKyMAeJDp2gkbz17wCb2wHZRJC49yiHoRtWdn9WtkY7mVLdvrqUiH
RsT2P1A2xrRNm6T/x4qjNDofShUzcuPbrCSn4pWxujSASLgmDusGshy6QAkPOVR0
YQ7qlPJEhafrgYOHy0VCG8Tmhh98FSNirvhSNDcFjI2JRBHiACtzF4TNGJ5HfqQs
zV/Ld4nqEgllZeDg/Wl6OCX3GjCeZLrSjNkunPZm+J0/sxVHJoJG3WGrAW/U63w/
o6FrDx30QfAFkF8SMiwTnbXgg49Ja+2NwJYdtxNOTZAhwgZxiYjIl1eXGXTiItWJ
SVKl0JXuNYWvWKEoDjaWYWYGqaX/jHEBMez4qV/vBhPmgSeZot2aN1TgbGaQMG4E
SHfsS8c3Zx8WAidGJpX4486LGfwLo9A1tdk7vUKZS5EaAzwyOJoxlywpZhc/hDU4
XLWZsLo8gPD4A3qT2bBofrBQE+XR+OSHJYDh4vvfeWvQe+xtWVq9vksI+LmYWVr0
HYU3GlbX0+y/SXn8YfyjI4fuCvdT2HJgRx7Tn2rd7fibfMGA311CbfZhUeCodM0S
6jvWb1uaRFIzllJCAjkNjDj3QTX9Um3cJYLTX60q1jt/PaovQiCmNTSofsYAe+gh
ba/v4XE6Adc1m4A1YXn+e2OTbfvBm4GYNoTKDgq/VWUnznnU4ZEdzbI01KVipktI
7ZtdekqiG0wBVjldHTgnxFUDZ2Y7NhkejRbiwST4YApJWgRdKeMzfRK/RTdbZIeL
RD0QuxbO/YsFpBoGeDgW2c6Zy3Ew46WZJf5QaNPtY+ZXVGFix2AoPSpjBwr96wtH
duPTA89lckLiQYaLsCACxOFdROS+HAB+htCi1/TCQtLQPc+7RTWLZM1l4RRmdyMw
cYcYhfbMd2BVmKk0aIqsN6+76Xd0JroP9aF45boEJx+XxyxEmbbrOXQ4ZrdeBqrD
1O/4dt06h/0a2DV8MqW/7F98Poj8sk7nFFRBRB585NCuZchVwgqimZ92ggm3oYkD
5ODXkjgbPT3GVqMdcGZlOrFWXRbJYvjYzuLbtoKnnKKJ/FZyHlhlwj8oinT5Q9+Z
DwGnMXZyq6Xz/dqjdsH1dUU9KB1tNnQEmt9vvG9j3twe2nSOoSL5CHOTiETK40ga
HXTuWPmxYqyMtaXjUmFmtwRmPMZqqy6seI98D7/EbI84s8+T+c9ZkPwTS1Bti35q
Bu1wYCGTj2LmMHcxGJIK3ItWXo/j2YVRPYyKeQtEhuBcUoV4JDX8iCybypmNYr+8
YasChhUYIrYBtp5cLd8y5C7/aEHeWr9H+WUIZBfES9XjfeC5yA/C1B1+9Y1VSuy/
GHen+D6dvB5OWv5fGAZnugN7pRma/XJqxT4yxyDX34HqZHtDx3FFXLpE6l9P+QjA
EN+TNil2iqigS9PlZg2ym0mVhZ1C2/NExceN2zA3KhA04bpWZ33SHwluoXEUZJsq
YF763kf4RFSd4c/6HLqaljrvXxiu3gr2vN2tKC0Y0/D6QJlpW4khE9V0tHK5Xuc9
1T2Dh4bGSu9OELYQ3+zx2sox9rlxg5doASEXDHup3e331Q1opv23ewBFFRdZmzKX
EpijjNoGQip+0rRGZgI3A2kD9UpwdvZCStF9rJer/02Xg8eCEHJw3RtYfHL/jEvH
diONiYKWCfhoA+1AW6B4orncDLq4dMpYXmtfokJPyrusMeGqv1uUMj1KDGyjgihr
khK8UgJT007hjiUQt3MStuJ/PosiQe3YyTl1RsPnjtpW1RP5/8D0D7Disc7B/td9
en/4x6hq/mzIpO/W+xydwtC99kzh+SDFSXb7tVqI6yFvwsW5AtmoPLBtNy012/BD
IFGRlBOrOct3ikFxAAIhAWScvTBGOKjxsptOUgU7jaSJkOid3iIA0NghwrO6mOcr
/BMsvxbGO63JXxWF/eiIvfPZchRBOzQVThYuEEDpskfPG+YovsvBtcZKbcj0boNn
TIdY/1EmqGCLexYqr5fCIPJz+cz+Mjja6wb1WqWN1lXHNoP33lBtPYIEI4Z5uYVW
8gFl8BeGO+FwUS9bFlS6K/e4zWLwyJWaw2YT2osbVMVgH4SYi/yKJPO92KM0BGOg
B5TE6Sd6YuSmoayx322Bl01v/lxAZaf7V37wwlhsCvu1tU+u0xE84Ndz4/ooRr37
z0g0ndUqxH0Ab9eocvb7s2N9jDhRfufi83DO4izY45pg65Cc48C2hjaBftjioy+8
RDbNWo2c7ax7tcx9T46/lHlzZi4HBzuFotZeTJQKj+EJPLoMalEIOljf5vhOmfNJ
z6sWBqefQTeU0ByfngbPnUWRIyUVkHh1ERHveOL+x18i229bZHPe2XIytsjTE+fX
DdGti4vVFpxMm6Zc0cQAC451+G696Z75ebQOUkhVM8Vb8UWMuqRyVvHRjshAHORM
FhlowdUugTnqhbEz6lheC/+Jn+o+tU+bGSQM5Dx7ichVkFK2G6InOdeZChtd9rEP
LUTxF4dfvieoyDXVjbm4+CJzMJt9G9R/8aTArm4yt/pE9n1h/WLuaigPiB0RWyLI
aakygEG4x4QBfUiQX249M/otZPLEn2ARFhSmWRTF3BmXQjjxDgwCJ3DuUSPzeCmz
jY/ZbRqglo4OZmvUJ/RRf+IvLriy6Pfz+3Kxc4Hy6Us07nsEFgcXTXiYLbS373ZN
xajv3xrjzp4pNtBXT0kXDzvt9W4H3i27EJBoIgXYlq9S0gs2c4mmNA/2SJbK7Yme
DkR8MPF1Gs76iEKVGW2VrkNo8lYGbGY6nZCb/atn6plfBZWpECU9qRa91nNmjpR3
iiTSLP46MA/TF/EXk8wiECP3E1yJ+HV9WELRDrtuemb+cfzuXZoqq4KAR2t8+hZJ
Q4yP0rGJhfeglyAoetq+tpVPjs6chZj6mMX2IX9WwRMA5lQqX5q0QXE5Koh9IOar
+80GEH6kI9I+5F5EZf3fY39zW23Yl9dB97JeLxtr1sfL/idXtHiuQGK6kc7HoAGF
Pwe73eq62qpHJHR4fd/dM1sPwDvqptYHOBpwb70qCb6ytU8SSQqF0FnVXvhOawjV
xwDjbKeXRtQabgeERluOOZtsmc7RUW53ApShxmKNQzLIvyM262ejADsoiR+Cis6Z
8V4TcguKS39b2lg6+ITGzleYQwqPzABRbaZDkvZMJ2Fv7E0Q+WobOa/Jdr+7NjU0
yAIWdviT4SbO+5gReY9lb5a3Vdn73qFJJf6N9vpVNcFoECKaHkTUgHh4Sh5svIpj
MGTlV+kByn0KFUMJqGa16pmCjsSFDl8u/gQ56hJl1qRqo4Yi1UtRsslYFvmPatTx
ntMCXY7Vx+BILiuowI9MlafemkGUkVIUS7J9Ht/sFDjiPvGm8CVfI5UtJLrlZ11I
eB9+bVndq1s+bjUNZpTtW4ZEGIr8qyKfeBr0riLExBOGRHWKT1yAo/vUOqvipgsp
EqOy+0AVKwFpCE+LT+a61snLtWCoPm1qGPbYBdrrn8unIKUYKGrkz3iDaUFJSJAM
lkhm4gYsJpnr6ZJlQwdgKmdjRHVjuWr0WDR5xvSP1yekxJtTw2cPGauaatLj8Mpb
bL/mKde1sFGe9wP2euqAmcZSCEx7EYmAIgzdZADTXL+pOyCstL6ANi3YmW+/o4mj
fITnuMq6n0Jl/L0kAhIj/4oiixOY8rMO2/9SA9hEV+Jh0QzOiUe0NPQXyZ7F0Sd+
fZKBsvgp5BbUoWD9Sgo4RjVQsrOvsvhhjJAXTQFQoG3OnAXdqrGKBArBbpG+PLEZ
YcEJkkQfreAXwwbZWAS0ySDcRjHF64ZESC6ktddj6oNsHDDcs2o5EVGAPuaqZjNc
HMppTZEltFt7bHgCbLnURvPkZi8/QLyi/i2zZdJoXNZEtr5kEazHpqZ3An2N6/Bz
AIJA03SduMryUptJFBugiXFr2rXHez3vYPqNnklvvKu1DygOSLzZPcEe02ZRF1qV
t8ar/sQIsJouB1OgC8N7Z9YGSXvoDRpws00IzHu7VIr+sCE3k9D9ZykYJflipR/M
k7vOtgXQ5VhV2WLYyem3B8u7uwUEUoxo1eg27eNdeA8tFO2mcKD36p2me88hWRq4
3GO7NEtt956CJcnLvh8lZgauy8tlEl95Hr7OSikEQEBpf23I3fsV7Tu8iDKqDInX
9Asj+hcTmRTKJncZlRMJeXVnU3yvCfTSk2K+H2Yi9UwiVovodlc3/I8tE+CbvJPJ
+HfMX6SQcCdRpQ1JxB7HLZmY5f4XsWEiTzbuJQghdcdecYBBRLsps3lMwMc9DcAB
8Mm/CDADdN3vVL7yppHRqeUO5Kwkbsao2e2E0FXYC4ppRNeKwx7QVk/XXrEfmrYP
1aVqvtlSObjn70Jmchv5l3F5sGE3qj1Vott1VZQHXTrFnI8fmwPdYpI6eal8dBDY
YvK6FQYjAjDBewwmfzXmYBttv8YsaXPfB/q5klr60FSePa+Wf0oMWRDBuv/pPIX9
18UofdmHHtPIqzuYeC0MBLtPLKykZLIX9AbQ2FaVmAgSq7TXY5c+XgpT4j3+rgfo
92a919W+Mq043ELu2ecBd1wIIQ7sMIi34ecCVp5vcK67s7aKgoxA7c5X/kAnFRsR
nZIvmTOh+wHo0RQAFEiZg3sAHzAgSK67oIsRZxppfofoSNf/Vcwky4nyMt0SqweZ
98iRvL3DhRS5o81sa6fCZftFY+x+hN/gG6mD0fFZeiDp6EmvRmNB/4s6tpFzQPYl
89LBbdDTWDwlAikHLQaKTl4JQG+nQU0w+TV90L6dPXIN5H20b2vLj8KrKjxDcUuR
8CXpPcDm9RjZfUq5/S6+hENY0DLk3waxF9bi7qPXTxsVxAJeYhZnBn9ygSOIcFGA
MYbffQjJ1tywrChG/sV5H1w8OFcW8jpztQ/iC/KNflzEgQkcRMnXl4XKX130i1OE
nk2S5jZrCy7aDUFrTbkcbOTXF0f26Bf+z5x4rJVCxGzNQqX6SXKp/E9SuQxzbQrf
slwdSEpL921t7Bg3LukbbshnSeJQNFbrujdCqrBryBC0yoLriq+gMMBYJbCLwEMO
IkLzCfWH3o0NEAn4BPcPmTgUK8p4dC4bdfs8vLZcq51ym2dDp0c30mmdt4e409U4
Bh86s50eE04ZXKk4mtDVdxrSA0JehDYoBkfYM9LjH1DHCgIAwvBHs29pSHmISrCr
RmtvQF8ODezB6qRj2iWGAK5u/YGLcseVwELR2XQu/KljfUUWH5Mx2Npg8J2A7dQf
aaeS96rGLu9DO93GH7b96BSkSNuxj0x+svgCZC7uXMFvv0p/ZZHWGqsfPi1r4X0a
+Di28pHNKGlBJAVecjGZipWSOckjt+AWvREo9TMprVvmMKbOefzt2JO9DKEgP0Xu
OHFvOAz53sgbZkfubJ6KRyvSNtALSK0kGJxUFEqwdAx2OcUpQt9oU1q8ZYp5UmrP
NTNjPmxYUl/rmfiSFvTvb0QEJX1dtRJVwjhLMHcVSFO0/+cfEfARFZk9TZXWxCj1
lDMjdyh0OWy/fg/YdXxAvTeb6m+NOHP6wvZjrtJQF96TgJdE+rfkZxjk/zAfV4qp
LOtDLZEqpGIeqcQmRZL20fv7R4kY6L9mRTX63/f4at6AoKHbtNrDnHRjzJCY8Cg1
keNIfmdvP9wq/0T20oxcFKAXLyUIhrppS/7zuvfcrGrEf5UCyYyO6vnIL/YGTF/T
a0bg/f3arvIeI9t6YQcr4AiLGxZTD1Kn1ipGlm36PtDTGv0RYx5MWp5w/8X4fAYR
MTzujdozWLI+Bso7fp5lfA8XX2IA8Ig1S9Xxq415xO96q4qXyskcFpgjf+D+uAnS
bwEyz3KvUFX0oyswzQZoPxQQS5vg65esyPnLrmrFdNMm2JRdbV39ZPOQ9mkfvakw
Iz6q+SYiiNZfKJNU/dMR74NGAvTacJn9SrPTFVYLs4qa4sXp9uW9FmqhYpg2d8JP
WHkXV2qWjn7/u/IcQ1coX8TJ1W/LmCWNRurkJlRWhv6rEVUXYm43mhTZNO07HPCh
IqfEr3jpGOueCSO1ALOXCMmL0Mawwo0hY7dJpx6eCusd2PFQpfcs+zS/RposDo6d
szql8KGo7zxS+S0EL87rGTpdK2p5O+6BWJBczMd9zlN8GJfSg3n5AOgqFOClDRP9
AC77TFvlREpulTgRAXjfNkJo+U1+rayJ8zI7LEj0IyyPcxH7BQbOQenL774SCngd
fz7HEli/8llUiqGPquOHRFe4bhZ5R40wzJBgFiSXT9QzjQuwI9o/8nvW1RajCeYg
v7HcVTNvCQgl/iQkVIdW4SC/jCM8QYFB+pAhYctAi8OhStE58FNxLaxjwDv72cgr
pf2NGrLjCoWHy7nNYpawQu9SnyW8XaJo6aqPt0CheejkAASGiTTAf6IBC6RYEAF9
W5DB2I9fTLVHedjRicc4VWA0zwaKAOxHC+sc9+97zgcwzWzESFeMgSh342yZ8AP6
BMx4n9Y0xwj4xxmRSNYba6yW0QUiE715w6TsiYTRDLFRyhacePJlAGk7M+2X8aAh
tsXqP9uSHUHtM06nYIRseNoQmleSMAavrv8HlZ+a6Mr1cBXnLcysc0OaDCYquxTe
F3NBaiD/dpU1q5PyAiDvLl8bGNURT/z4ZR3oymmuXrBk3WVczl+TaF4jC4bwLquU
YP5dzHP8Uz9BJGg0y6zLWkBRRc4Pv0HZaDexdNO+L+2RDz9w/9PL8Uty4C2/0B72
r2C+ZN4OF+l7mrWq4iBVaMY2Z+wVC7/VSp757ZQ9syzD2TT4L96M231rd8g4LS+G
bQkM4I4UPXKiXSfRx3AtRXYuaBB6cB6AYclVFj1UJD99fbEsi2A081Y8fKfIagVX
FQek9hQ8xtqJwZheBnWKN0fjtF2xtarL6aH6Dz4o7xrCiz6gU13XRoe54yj1JUGz
tpUBLgdj0XQqiieUM3C+mjN1AwcpULNVK63bfUdfSjc9bevw2u6S0Vr3rB8QjdNr
gWfkcP0xwPRNZ5jNc8M2abxw+0Hj3Q/sfBQLzMqgfmvT8WalYgU1hOmUcsDrL60J
afIMyppTAQE/KfsDaFtfy+OeWoRFd9qT6Zf435qPTd5DyENZ9lE/sMpTFq6/ePhA
w1aYgPLVJbwBGnR4HsaVtwC9Yua/q9g+TJA7RuKj6Qq+Dlo+NhPHAHqsGARV/JbX
OkGFfSjEQJqsALsKM1zRVZyhM+sPOZgVGK3/GP4rCnpltk2sRpKKg2wrjzQPVfZR
2x/1oGDHekWBvnW8F//PBG8XOEHZEE+67NF/aBK6Ka+vO+UY5NEJog3HWePncZac
5qF7SFjBOhjInHcDC0o/Cg+kpGGamRmtQLzA0g9FtkyxM0CcVxlDsaPvQ75UaLI5
03Nv5MqIHoAkQGsaJJ0pGNv7pJcisv8s1D8w5V38spABFnfXBp6cgb/5H1/ZLEWx
olZZh7KRztew5FVlOyyJXWVRMD9I58y3SYV28fl/VsNhYfr35ih+P+4JCzTKfk+q
FmijSztToHkqhj6tbBrS2gRda0HGJZtQflt+j2I8SqatncmIlwC3g4wSN3QLMG6Z
f7rGg0c7CHB5Df9/sTxOHtr+SacDJIUeHd6skR7sweS1w1yaZjGTJwfFlMg5J7Rv
byHpYP58v3RP9TE9spL9Gkh53TOZP8omJA7MYsv771/EbB8mrw8ASepfhnZZSO/k
yPuognSAJuHJr5y9ViCwJgu8JBAS2+VBey0BtWktWv/Ckd5vb0HBFHW+z40mIF6t
VPPUsBUisqeSaNzZEKSZ3zJ7zk7wRxc0Ce/BnvEJb2RfwZr9OIMnrbNOBE9wyFlL
2FUPgfZ5VyUGh8rKNASbRtz76+ufyB7dlVk0IopnWKbF8f6xv/CwJgYFAVdaBaJz
ShjWbBbvjwslcA3XPHPcqpYVS+Vt97KsQsp64r6rABfE/9gErgVvPdwiJTps+Ril
kfetZxcyL9ygRcNA5xKGCaiwFD3H1RyBYe5lEnvCjbQ025iecMKpGtnoGTIl2avb
vLyNBIWaNKuCcDiqwbajUljct9pBuQBQoKAb+qJ1GVaQR8jI67IL0l/QACsF4mWx
g9pBUINGRbN2zuPh25JjAyZe+Oe1xDgey3jjY6/vNBph3SU8Th18jIo+0xGA/Yg6
hBZ9kmjz5rCH6ob8iV7YoccTS465pVDjRsnj6J0LJ+zvQmNmDtVDD4+RP4O56fmM
ITM88wmM7GMVCICeR7oYmTqriJsx0f+PXI+HoOLSt5G7PYI/DyIFOgiyNZvLHN0m
/pVi0VZCkYfJQABE3Cm/yYakl7CKC7Po0vLFTIuJWld+6fyBgqHhtp/zQGEdE6OP
MacjAHJmlpr05oyCvxvDfB5tbP5zoVNB5QETZNJ++1RSloMzOzmHuEByibTo416L
IPU6nrhNWrsg4D94hrFqhoTasKEUNOjvByeBhBj51Z79scO79pnapeu7uQlvCzig
r/kADi6JhpZPyqKjNSoeQO2wjcIPjJZ4IZE26guloLyllvFCKWzxQvoAPCZZdyOD
92S1fSMJvMOSAJoH1LKXKnuYt7aSQxZDkDwiRSsAFS3T5sKUKy2zN6DBnIY/ldzq
OgIairX6ZcxY2q7RB75vdu85XMyl2VzXKEzexDpnp6N7R8esvh6eMq+fgYCJNHKi
G0Pub/fN/L31XFittRvk9WDwlo7i0xDQcU8kfBUAuyLaBh2d+JbDlHhVdSeaJ2n/
GXf7phuLg3hVTP6d57K8P5ml+QJGBEZeD9BQw3jAdI6aSvDaMZPkgJRURE3nTHv5
GirsOp49en/wzGhQeWxEJKxBmKWD14s3jyn8Kl/wTfODq2cvt5w9coiIqJ6H7sgt
i9XPx8QyhnHYRILv4vJDnrxVmiH5d9uAjPjTWMyLDP3xpElYt3MmuXruhhAMd1zm
tABlTb7mKhJUmfFAiu9uloliRJDaYAg6PCO6br/itk2JopMiFGqH+sZsyA064IJF
TWtZw4xFgSSyIh6MtbFIt2jnoUIWUVWy5VxjFq3JZgbvld7OleU2fAgfkt7wYekI
OUa6QJRRKZnqvZcDVnif+E9ZL90AZDChsIOymqN/sRoW7Dd//Cl2hm0W/HlM7jC8
NhKR1164SWAkX0yiGfF6ZrSHojGgVHsezw1zTALD3lkdCJTclMDA1KtLmgh//x1E
uWBVMXSGqTMX5G//+9axDlU7EAySaqUvVXsK0oN6twoZBKaDjU7m0oPuUF8xZrM2
uQUtgfj7q0rT09plDOwBDkTyIKw2uJfKlukGqTb+oSCuNyC/Jw91NC0wu1v/U+yO
x+Zb4Pim9kX/i/YaRCYJ/317flRu2rrfMDfj5p/W7Zzl+WW1uBCNTjDlNWZRVYsZ
2OsUtYKVh9W3ca9xIqhjmGGR69T+O+29SFAHd8NjI9RSIBfPl3+6/Ql/0cSQQFjx
EAxTO3Po+v9Bzs+f1UgEuazvwqfKGSsKx/5dusUxwMWwPNFvl5v9h6caGLWnF1Ah
ef+/iVlC6a82QzyD+X0PpLBbrgZcevm1qM9P8tDyNAYLMZymgZWh0GRmJg4GzxWP
nD3wuf5cM/rPE2VdVhydlIn+0QwwQtmQn3Pp3KexUg5E7e3aceVFyc0eByWaEwYS
iSOl9R2nPNJSRS8cXcXUvswRn6qg3/+g7Oizw3lz2j6Y1W75m/uZpeUB537Rrke/
PuGY7qDIJkDBZ/FvDBCdyo0ifpYMZsB01NUwo5HimyFNlnVYS8Ox0P3eppZcpHgy
6EKuBmVEviUEbvsHoqI6EOqHM0y1F/JPzVwdOEp63gV61zJvd1vjbj0cLK5LKzGs
GwP72ieortocDd6CcTCHvIrTtVHpbSC/NlSWxfCHpslQMKvuUb6/tfkYHkPSalLh
NtCeFxzmfDMeEmOnH/0wP6IcEQVia+gZGeMC9z6DfTzoGIFTLOc4Z/dl5MlzIjon
0b9tia0ktGe9KZHucAaAKyu6t5n0tJAO71+bjMEhVxoZelLVyPnviVxqN+Ut34OD
IrxNtBTXgk98dXvj/p3wllAlfrq5W9zv8+7cyPxbY6pKgCLDxTjpa7etIScpcuOE
DeG6fJS6O9X5z8ulDSzEtt2u2/BfzjV/aam6wbB9okZrl91xMuetu6JZ2M5XSWNp
n4cEq/ak+4aSZegb3LmOHb4Hl9odK2O9LfettZVg1D4=
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
I5dIKknrZJM0YM8FKbiVmktAamm6kqAJoAprvm0HyX6bFFHNl08RXJTArrt+I3mc
mwg03RaMxkd/Nurg0r++90iIp+t4eSvckpEGYmpgDbpsvIOSm6hasubEM1C7PVFE
3tcozPA0mzU2N+Y/7TQRRcr75ft35JItxmko9EE/6hd7mb2C8a7NreZpIrv+Bpi3
k0ce13L3iDgxvvfhMwCk1nZw2O3ddCly/48EgkpgnP1F3DokZK0r2lxmotKInL+q
KLfNt7as6OkokTAhCk1M/6n/rwTTQNHqxgDVhVlMVlVIptphSnBOaD5L4gHm1EP8
18r7iS6tgEQZ70nqwYP+TA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 656 )
`pragma protect data_block
y79novoTKB6QoLexNzRNrZ9lL9tEGWrxiJYWctqfexRlSf83lk8TvR+Bp9+qe712
nxf+c4eKMJdxUP7cMFeT9vxwH+l8TenlOtU5JekefnuqahJkFTvR9fZKzIQqnSPB
//o06gKBkRfsLid+6WCE0hubUQBbZV2TDqxsmFVQ6TY9URkdqfaGOt4mofFDoJxw
uzZzwlGS+ginkfZK/naVPexDd+QuotLgIi7xPjBLK5oPPmemEXdISbfAwyhCCVUm
0MvbRYmQdMbT39fN1eRRUc8sM8kGhtBIqJJ5eqEF9igjIP0k2sKmhQJesH1eFtKM
+5LmSBAJgFz1GSSk8io0Nvliui9Abse68ZbLdTlwrUAhSacdUtV8ZX9NIijuUOK0
LPijbfxr6tk8EVnC9bHwrruViqjUsnWVdPX4dSLBZpjuPIOO1qijbQ3o0kqOVvP6
rc58tCq62j4AVbXahgbLVWR12llnrsnIlgDjrqecn5Iczag241pVBLpp/3qZ5L9r
gXEGfys4K1/O5B4T0Hgw8CR6H13/UZsQII6urgJ+NnyvuJ3fcMpBbTsyMRKTgFBv
dDjsN6EBTp+W8EiM9oBK+AZFsydEYQzAeBP8OnlFklYVcGN66Qou7q18S/HmGN2g
ehV+nYkzGE46R7olIRyIznTM2oZvBU/PUMgzGRW19vGm/u/g99XUsTA3877gtCQb
ikrO+pUd21lpfCBuv3afj+YgDsfvm1/+eolMB6MsgTHyZ3P3p2+cqUPb9FV4j8xa
DNOOzLjYWLvhDzRSsbuim+LMujUUPowVy9+S7pPNbVmipJ6lQO2Q+nyasIQw8U7K
nVvwrbrVRVuIu51SPOhZdy39eCp7maycQeJgL3uzFIs=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
arz9S3q7OpnbrFiJlItNhY6Bv53peG9zlTftqZMNSPzyLPgy8KAPY75gTYghTYdH
8Gv4jC9B6s8quJ7iz6XbBskm9h4pXZWUulETmTkqZE/NhIcuXA4bMqvYUwUdVAjG
4oP0N4Z7RPLzAj4VutjJ7jJPmDgk5pmP5nTt9ECjbuDBIGDC7jufz0HVAtOL2fPB
psp0O0qkNUJ2FSNVJJkUaj3ZVEwCOUXKOoW1U5+Jp/8O6H7dJQZcNCTLthDvEEnm
WFoBERBrlBLlmkwS4wibdV3HdiuIfUOvQ+KOKRB0dFgwWEbuh9HTUQgkdw3x4T7r
+nsKcbALySl6fYQj0h+g7A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 13024 )
`pragma protect data_block
hSm6uP06ZrRWgMqChYpHhjE7zrFwZHOL0tQkaYv0YAcl1x+H+Jtp8Ff+Sv8//Le9
K10I5A6P947zRNEEsJv0/pWuePH1UuRDUKbl7FK4GhuTESU24NEqIqkhAsp8LFZB
vrdrXS0ujAL7u5Ffq1eyVOM1o3Quhu9cZRVXfevtiZg3s9j/6z8MnZi8vBAMxG8/
IFizsGEdYxfY72xXjHyCJmeyiw7qSaHLGTf+9GDLeIouPcDK0s3JxCeSTglV/t9z
VCc6G7oMUXDMZ5nZ86NWZc5Jve387c6hdT1GXfpNQEHjTK3VVi6q9jOdNdQTTm9S
zBnhsv7HN4EyPwdImfqa6/K1uVf/RKdMDmXNJX4tDwMZLjSFWxE4m4o2Cj/8TVIx
s2FPTl30hpIY4ke9XwBtQPAFvED5Qk/2+eVL4nWKVj3VxV21hBCapxNIgd6OcSm3
vb24vk726gBWj6wCyqEDdMnmmFSKHYeSSTxfhwwa15kQ0zzbkz65oWeWvt/lbiRT
7JSQgusLrSpIzI1ujKVUahldfnmDeiFZU6Bwi97JELDo85VfMlm4tmuSviI0ry0S
S8juJaLEQl9m2trBFbBCSKTsvAsKC9Ze3LzriSURAbAdEmX9SlRZ8oD7tLvsofK0
Cv4K2RBbugEUgYFcmBRhyAH2DtTKzsfIX6ClA2ZashWVjnWlzF5GSEJDTawCsfql
6AdYFR23S4XmdhoM9ugqdg/4U6lsCADp56qiZjbWA4KaL1HPeg6Xlon8wyjCOogx
/OPUsjv9s5ERYEz00XWu8kV6Cd2DT5qQYR7XviNsMUIKQG+RbNBsc6M28WAgUXup
XCMc8A6KUPK1xZP3sF9mbfNtR3Zu342WIMen2VS9nmROXEEvIXhcM/h1pKDwt4tz
aSHm+No2lATEFkGVLVWHrlbgw7mt6om1OuThJaZNVT8YHva9HEK03Z3Ubkwi770C
pNOFY8b7oRC5xugugp3Kp7YGbie/41+i05Pc/KHsflW+XeM59vdrIiu23aYQXQAd
kll1hxbmouqfpF47r4b4bAJJCKMa2g3k5hvx/oyrWOR/pF0cUhlHnYgir70ajXxX
lz79zShGtTgUcC+nr0EnUGOjT7OAjuPSAauECGLaDKxT/7Ed30x7HY+si6SuHk2Y
WpSr03I9eTXdNnln8/tWTb+BRKzU8Bh2ejv7tVuOTOJURmRLJXipURW8zjkBRaSa
IwDHBxlC/TfAygpvhCCWkpK9orJuzLaXedsRrKbXoP45hcRW9wlyB+Sa+LbvJ3NR
bMR9vc317eJfkGO664KcRe7N5QYY0gDXsK4q4nnQfuca7594B8enjLiR+VCIICZP
N4DVtQI+D1+ird4Nk9Q7UxyjZlDcYBKxUNo6c97NWV4D+CPwJHHWjl+DVpK5RH9i
QGOCtXSC0jJSrGJySG0dW1vp+ZL0gShaQjswqmEs7HUxk/79L7PRQlu7yYCvsyuW
nzxEW+481an2WbBlJb0K4M2saP2+R55L3xt0umN2uaXnNvT3/WwK5nNxdxMXsCy5
lwbpzplWprWMUD7f3X4yL0n/m7HVuLWeAi6WkhMbYd9KwgyY3SnUbxkJREHHQlmV
gCU0uX6V+9oKe/WZi7lIzWfc1l5rFtviiX+cPC1s8VJ2qgZveMG2UjOM9TEh/VZt
oCyYc3zi+bpgVwmwTQYhoNER70RwtE8jffL/sFRNQQuStQvbqBqQDHk8LNlzjS0H
OIg7H72OsOFyb4i97sFXlgpohStN/v6I6jZQKSB70a5MFXyJf0fc1oWKVjl51ObH
JxNVZtiS09x/aE7Q2Lteukvz+YFGsCXNVJad9hLT/auGIkiB7xztuji5Uggg0zBo
zG/iXDRYteUIAtmByIX8nTl55yVuwwWex1SnG6D/r7cQvh1AS9QltQizMG8/qsyl
+3YNxs9HsBR1XymjIBsO+0b6YWSycG/CasWrAqA6PI93uT5zMI/pdrxKktGP5bth
eH7VZdNTAxvHnT6yJaJduISmo8M6WBfQMi4yf6iJZQTOF3ScjO16jj/z0QYtwmfH
qmOELn/ReQEN3SxeoFH6zPK11prI3mjR0QtCo5oiLNyXozPmDzPDJUwxnpdp2o3u
+R6/6t7NGpil0ZMLIlolmWuw6I9ZfNYzr88D/+TVQHTQFAkIqkkcymdLZLJecPFy
I8Ae5tWvqE/V2UFN2mTNhc2vTB1wm6VF3bg1jCFmPu5PbdT1Hl9SMT5EctJ69wny
Fziu9O+Q47ODLu8Lf9+0pk6MXPcG3L37FRlWgwbb4/pIyUgxxm2BB9Hbs/v5sEF5
Alz+4Zz8KIEuEb/lOeEDKan2GPK34hNudtzhnLTEr8/66kJmI87CfCBBZHuIueCh
p0I2yik7LSaDVy0p6PvlYbyOMoROt4HG1Peyr7QGkZc0Ttf6s8QNujZ3O4y+bEoO
NhICLxQgVYb67Vh585ulvIgoyqMLtiaCf2dDTgMP5opHzU70iqNXQsDDSdUIEQwJ
iODKlF0yV4yCyX2CQVgoAzC4Ld6eh+dw55uR8HuG65cVhUUyPNjPPMEe554u9MyV
p3QCZ2Vikhb85ASzppROzQItxECvjZvLxRoJL6rdJGEcJLMPjpP/zVXI+5PyGFux
kmvlqvhGMA+gagaYP4q/5W2pytlkrRhSapqVqY1swc65y87NrvUN21BYHlGw3Qzy
T38U852rx/9/aqV+f/O75IUYkA13dUJrtF2XWxy2R7qaFVkrTISfwvFGKIpaAE8i
nxoMR87FePSIz1P6QRa8fAjcDiMn0W6fuVNdOUStWtaW+fX1zH8TjawsFtXyLCBE
GMPDsnikZJFBKx6nH3uAGPI3+th4S8ZlmQfXtIUHFHrZJsCnYTc1b2gjXLSkDCOv
2DDJWyotKF6ubAAHm1Wu/UUtDIkmU9tWGCOKjdC6cXkTwVQtBk6hiUOjaLnTucMi
FtKbB9Bh92MwQ91U/0WZvrO6GvesbPyl0+dh0Ef1sQuq0QOoHpuHoFEakhe2PRPC
yf0zp5VIrfx0M0QuoyanYhYZGxTUXBsjrnmzlvcmoS6Y/RJJ5rBdnj1jSWx4BPLY
NJs5QhY+dyceyHajJF2+RZEQJxgdjhb+o1Hee9mnF9gHzpYGYQfk0wYqG4yCZSZx
z+r20sKVhLVNK10kNq/XWeX7lbCz9xlEbLyS8eANZdq0H1q8B35xJwvcYen4Tlph
+sey4OsZQkUaX1WLyrB0IIWQfw+bGx3bVShyXtiwEx2pz3sI4vSlJcP2AUAAjftZ
DHoEWT01LV97dtp97pUEKrYOijwC/Fn0KDrbXI6PnDWKuc6tBWrI3guvrIF8h5fO
jy5JX0GNqEd7wVHYo1t3An79L0K81tYXHVx7rAOiuk1A2/JdxScEqXonhZrM8sO5
uStlvHEWx/XUkhkwkjpFuELCE7t9eAYnWwLX+WZK958xeBvI2ObU4lDDzVD87kcn
QpBFWJU2mum9qxrEF6Lr7QK0gh+Qw30kLx+qAw1sInUaJGSTEVFcy/jfFELueExg
of7sMvyHOn0krDXPZ6A/pXemfNmsHsSH9Qug6QLVJVUNZscz3/b6xiaX8k6eQAVa
JT5dEg9PkNVtkhfOLrQ/puEdYVA4wBrX88N/z4kWxJ7m4xalCmWhPQkQf/8BdBEo
4SMQS0bZKB9utBoiq1DjpABYIpjiveQLf36pXfAgz7pr7iGYrYZh/cP14FZ16UVQ
Nd2lnsJb3i6Rg7uXSqzqrSh6RgVGRneYV22nl0nohuWWU7uFPJmmlIH8+ITFt0sQ
mYWsw4FNduMapy0aaLCiTWK1IGBFLzhVkxOj2ORokN7tI0/fNRol+AkXx4vOiui/
k4zUYWgRRY7a/mQZg7TPma93Ps6rwO7X516H75J/MaCiFNHJ6D/vcYYlsZtBi4QT
BITxp6Hg71HUKDWpcf6smEbummmwj9JT9i7PN/Wtc/u4ZG5xR5IFH3kpArNzN1te
PYW6TMVCUV8WtHLfnYfr1wcnZIu7HurrtNODJVPBwtwJQ+LzEzF6wqMTxcwRbnWk
AI8gRA8naH6ja5VwEZd9+Dx8sNYsbIFjEVDiM80Ky/eEw76X7P7PHOZAHRNJOkE/
qwNWfilJO1kRgHg5ftrlKkTn8TKILWzb00CQd9XWO+njB1c8hXB+EKVBLKZTp2gh
ocHHgVAu9rAqf6oFl1AUHPDKhSU4CGTruI48r/SGsY//fpxgfD5RRTtGrcTz2vmO
KD8GaaPC8YmXhsN4fWQhsspjULzsNlSPzT0P5mB+GuYH+5H95dYvCW+FppZ1Oqpg
JLl9OEvp/jwY6nlB+FEXzZZN4SWmdy2PTYT1cbOdUSmPsuFUjSz+/y0qBpjEmMIH
TFuLWHLUP3ttrx9AGsOGQwf78UTnSsVfual9GgHqeOmYum8Czd79hlomigNbs3Ee
/wmECY97viu1it8U8EhPk0dxNI/xg73gTV0JPbNyaCbqQDkBe0z+o4cs+3fH8X4h
p4dEttRMSpfn8neDqXTN2vXIOPYcTGyr12ZuKa32hfpWPM2iPovu3zdyDNERkXTk
M7d2VsRXBrVwHNWKVPIgHhqDGSsxtWlubl0PvbbW1OZnFxUmLqPbhc42Ytmbw45E
U6r/ESy/iTofISVRJWeolrJ+75IielivHNufPJC30TVkwMZdzPYnTXvPmGEdwOug
dWdJ0EecxWDv6pOz/MpPPAiPj48u1BCAq0Sy+2CETYxFjUgTSA/NUKd6+Y83JfVF
EpjQC5tTkp7+ByXBvT0H1hToorn9Ns8hGdqly+TOeccsQibTw4AlLPsLsIHio7x+
adXXlW83vOEHSSe6FVmasaz2Ha9ioqfgDVu4LBqmfFDrCXZcBSR3zDNbc7h1ARIK
MxuetL6TwatQJ8cbgrfIyUeC39ex0dnR7LstqTBzMkhWxfjzlJsr5jdEoM6OCRJA
38bEaIEP2Y0JQV9WyhSEkXr1ZNCokkOA0N1u8iblCiE2SFD+ftXiqw8Dep42eWrx
6GH0NFmW35QCBvXHztVp277KSgN+w8Ob5Lzp8a6aLQQxfDwfLYH4g1dqrt//8IS+
368bPd3+kIkf8PQw5a+VzaVJzfkwQWt7u4YBRajA/+2N/oyof9GiO3tIqKeNXyRU
AVQ9W+9ykhvDlg8i2XnW0mlFKvwos0AD6Hpb+z1/oEX6VYBW988d8p6kzatXhlZr
pD/jOUSfAHuhInP7Plz396qrKrliG/Ekw5tEFy9vmKG+edh3SN3FomHntsXLUd3v
UfT266HtNr6WLZ/hGBtSGOp0YvcLd1IUR+WYjV03Ac+pg6OV4Xg9rptwqFiA7Y+5
TGbNBQoMTLp64tC8tlgQf7AlvieWYfnK8FXSsIU4KRabjdGl2Z5SAdZOh+e/3hyt
KN86rGud+BQAa7qRA2zCcqr3Auc6EZT79+5X9zpPV4L0uOtN79OhM4G1lQuro55G
n1pvnguEj7o+PuGeCYzw8wgLpXEihxOg6TCE3gR77+r4eBypn34cXnyGKkQIedqG
wXkq6zJ5qZypWyJDviRaOxukvW9e/fB/IGcncKSCDxTMtZawOhgSv5xlVSFxjLbw
o/FgXYk1vfAi9zctVpEA7PfzZYZgCpJqYaS3CR7nhn+KdYMAib5IdHn2lYb5dDP+
aVJppd8dmONeyR+U9OTYpLiW6Up/yCsfQa+mqOkEA0dt9ZdpS3zIf47KbZfJ6r6h
0/FWt5GJDyj5NX45wgKTYfDRGITWVX9lbnzto4l6uNeRIit/LSdMfisZSzvjGV8u
1PHNy701hbF0ynHozRnAGyGEwgAbUzFRoUgYAwsXg/h1e/ZhjI9/aLMbUJysgw5g
YrDPgC3ROd6dgl08i7/aNQHLTUjJiW92RcQ5aBg1EQCH1qA+s2XcC29hrHX0FF/G
wJBsI9qV4+yo99fwo9M2PTr7hpR+mrqKowf/wgKpA0cNIRHaPQP8dpdHoLmq5xWP
F6cRY9PIe9EqIe5kS0kSSoCzInAepme0CorchJo8UO7aCd+Hu9tg7zWjqq9/7Vle
/HsO8gICt0ZiZml6MojynB0DUW1d3PRKYBuAY04J/ScKJLYlegTQbTiz6dZPn0iH
sL98RxOux2UsqFvAImSwEOgnvi81nB+gSTZCSDbLBxw8PnQtNTQ8y34uiy7Iwcz3
DRUqLXj1BLO6fbMw4541XwHvvtHQGV7HYcFBYfTltJlZpH7xVZz5m/myE3hOgvzf
/DvMW2QVfxGZRTuylfotA7S+2KC3K+FHD+E+Fk3E6vmWcmN5dbCz5CevQZBLAH4R
jiY3KLs25ZKU+vZfyr7reIJ+bQgMV6xlfATpzE9djeWp1SyP88zV4ANT42UiQ2rj
3VxvPoG+VkEcc5nP3Heu1CbupPdWf+bDm6jFdn50Kxhs09erO1km3I0H/ACe86Pf
sjeTt0zh23X6YYXeZhCNtHMoZ0q5FLKdsSVPVW1wyeQt21IX8aAcQFGjyKQ8Qr0d
jGhn+ziFQbpxHWlh9dsevWmn1aaQGXWLPS6AVeQzG0RNXhD0rw86OBO/SzynAf+4
D2WitG+M2QUeuAex0r46fyTbBGt1CdUytpK2H1uuk6OMBsLR2pNT54M9vVU3zLyQ
82WHW9JfTSPD0nkLZ1C0BpB7WsPLIKvM4i/SygG6QP2Xa/976xfBPdDymITAIb3V
l+k4y0g6uFAjAfJL3g+79i/xvK+WzLEfI4bVX00sZf2ry0RmE6oqX3dutHNyA2P1
mcIczFbbGa13TicDAED7H6nUmiYk8gkySF8cZ37uIgrqjDgY1Puhd1VD23rEDnjc
FvPQafc2v/QllbK3dAfsfjt25mjOm+d2q5QBqQdM+oYrHm85jHA2qYFd6fjBF7fn
9zNY3piHyA1Crh7KjtuPkFZ2PVDggk4wy4XZtaT9W/hZRRowCBn5hZUnWEHVBCve
VkqX/1ftGtXFWOuHA2St9lIMAVfP6LnbrEddkcTcjjrFvd+6dvhqQ5a1NI84FFGV
GJucRARVmxYdJElUMR6GnOsJdH+OO0Vj1wSA2mcaPvUgiarZ4RkE9vpXHSx8XjPq
WKRI5yaD6/Pb4u97PYkImBYcNVLUW4ZdV+yaF6K3r1T2m5mW+PHjP/+lwBp6znDG
71O67Q4yWMLrntaxdHafugNuME2bhdWvuMJkLqwAfZuIw7+310p+CbCM+xtMOxUC
Ghn369zD4xE6XMvzcNQWT4OHyJefRx+aGX1mo5WZ4bsMIvifKRdbJqxN3NUTGXue
0U5qYUFyD+fvzc5lwqJRTLPvJwkH8aJjsYcEXdGoNHw28zRoWLYBiZvNtXTIV+l+
ru6feHO/6NvwTXPYWaTP4WJmk/paHkhCGoUOb1KP/JZ0XOquovt75ClaINveN5pd
OqTfQPusTVuaDeEwuh3bzX2/CIJlODGYCk7pC7PrQDdlWwAdcTVCbheGbo6U8cn5
ByuqKeZREJKggy5fYzyLdUh7EzhZ+ftf5J5WguupqWdKKLu2TGbHWhYcnpEh4YZo
bIwGA0fNP8tBivduveg/0EAaaoDCJ6kKMHKnuIjVa7osNHlsuVq7MrvZA8Qr0MNu
50TVdiXANPwERRReYvJvDmED4GPnv59ZB03ZkUw8KcyglZNFTemViWPBEL0rbAxk
EctpDQbBojQ172wNFg21lUEb2gMvP/k0212cwOFWyUTOxchvAwYJdjZdHJvJrInp
7flRoeyGSs/t6ExFkCnghK2pnCsbNbYlNgrpNTJhPU/CsNLqI1aopPI4D5AgVCpp
D5qguS2z5v8V6twaag7Uddv38nToiqwHzADNFQ4r4fMpVJBGz1GGrd/wFe0B1iPT
PvX1oZaD8L9NcHNFXCCFPuUadnd8HvWZf13/oxPCQphLHxjQRnSOk9kgb8+CLmLf
8hIIkysXxDKMR6RkO8Hmkq7GqhNyDJR1mEJcYGhLlDX2RBM5xJ4wF4tn9HaSlBcV
auD8gRtQLRcSqQVBUPQyxkJCFlXyMhbM59O2VJODoA3nKq3ETuT39U0JDdicRa0H
aYvLR0ZObJDHWHo6RkcCtTxmmCKwT5RowJcf8ri9GPFW5BPAYBkhuwvruOqMFAvL
QyJFWBCK0zvrMQlczVmZ5BKGPhZadtOiXur+zY+kRqtvyR4ShrJM9405D4/P5RJ5
tuHie/UJKk4lYMcDzSoVQVTIElvFeouASzh8ATq1CRCpGk6aR5ldu5UHfA1l25sM
tQg+hWWuEIpto9ULwZywJ9Izf3KKebrxQtdUXj17TREzami0hhdDEwbbpxJwV3c9
LkJLbX4Z8o9UMRor3iPZyLkNVq7ekKTOzmwocBGvUJZVhAF789iYf+TaMXjIVyxX
oz7Rj7OCSiRYoenO2PGXGxCBwL57lKIK7pwrurA9vZeRzNTjS7JyvbKGr2SdzelC
5EQU73+uApXkKhz9H98q5fZ3sUCylEFd0LxZmmj22kG/LAcEPAaEglQUtbdrPlOc
+/W67LHMJURvbNNgfV2d9RaFaaw1Jxwf7VA/Tgd4A7rKcuO1mNZYjwfTODGhZxgB
FINjYwriGox/DiOhuhquvabVcKtXsDdLmMdjgGI9Z703r/X2GofziAl6aVr7Pq1K
yPhac2DMha1C7982EGOijEgQJ9Aex6MAl4fiCnM/fQjUaNiCAaM9LaY3gO+H2Me9
Kh7oGZaeGhNaEdqnLFBKM02Z5XPUfHyCX8tDFLDh8EphNMAc4Rgm9586WUeIEtR6
YZQKY79HIJbCNc43hObVqWywPHaKpo6D8jL+7DWYez4cY5m3mGnCgWaCh0bLB0gV
NttSDsZum6E3Vlx2hiRk85Mn7z1Yh4Zd9qGzDnmgL9YQ6lVZOIG0cRoBf234NoQh
SANX0OvxoqfCTZ8OUDJXWrKFoC33se4qZqg8mI/ej3deAjeuRg5yI/htZd12S9xw
3wZ59RKNmofG+3ljD99V2/hIp2cYNgTtjYXHmJIcWmKtU5b4IDdmF+KdLNuv8QN3
WKLCIEY6aviLFILdIlP5iYMmpJaG9IXhAuljVf0Dgmc+MJTeJdCak56mdJvdM/LR
x6GQFbDHSWVWDJB1CLCSHe5rY41cnGUTaUt+vu8p0/sTZCf4nDLM71ciqHsqmmeb
5OqSEOVudW9cXDieOIlH5IWgonErJROV1YeCEPQd7RYvSYDgqcP3k3YozT8XhoKS
jh/YGS8k8o0QOD7n5HyhSk8O2Gy3dTF7kcuNNZX3hEfYDILiDVcCIboat1YJfjkf
mMyeQpa48GFc+BLf2OeqWMuIRudyqEmrzc/urA40ou//gSrubxsR0wNHpuhkRoa3
nxw6hkgNyPG9QpItGKqn9fqmFAmwcXICFqbqzLyWpeK2WzNiq+YICdvb19f0pvoC
6mPlxDj7Kc4LPmwUQSm6LOqFWt7P35RMjQPItMWWOAUoMaj4eL0shbgU46ao3/7q
woaTFz1HqCQNI7ewdPmmI+jqasDfD6zmj0HgHnpo5Qv5lp/LjIfdFk/FOc4dgPan
ZanMD/pwRy9yKHmNFzZn80hMZd14GIr6Di4hPSBWurIezKPuq2o4+WBAa/ZlgjD/
q+tMzY3VhAmvKtBEkIMDGO7UJgWcLjL+X7w4BHvdptHBWJ5cjEG8feeH+7espLpa
vpjRsfKv96zoowe2Lck9vxB9kDumClCahaarC1HdIs7qQJzGfr62f1//ph4PTbDy
gkkrdPI7AMbaAvsxMwYRZT0ubTykcOT1tCI6Z3TWCvTWccQ6UVDyO9ood7/TklTP
ImAuvh6TIsoNA8ocDhTFB9LCerSl3X2j8JjuvS1T/2AzwcmTHLw7xUXcqWMzBGSf
I6ACfo4XNRmXXPAuomlwte3yERVK0iGY9pPEojSpUOqvLRA+nT6Z4FoWpjs16h1G
18j5UJto/pQbxP99cNeYSPg+6pq0rIw8syRZDFOUxuKSwx70V1MY2FyGMEgfKLLq
TGtnHjRuC3pS9Ebe1WoJG2vnXPx0I8en2YZN5NW61vgFIJIAPSENgzOucElq2qJb
1A5YLVFGmmpSbIDX1/FLoKDa07qeB/xPhmDkmyF3mBqV+tEvB4Nf76MQ3OYziOcI
B5Jy8J9vbXORKVy/469lXDUg2PjuQmdxLZy3MBg6bpMs+0P09rCDryXCMBLBe5Md
c5cz9wNdl6QvMv03cM6AglGa9cmQtxN04wr40Cl8ECUaE0Ttx/XV/vUdcq71BA1i
HjVskm066j4OYTupmKf0VKZq3qQkQkKcJeyRLqK4aSQmw8Y1oDZiLGFBrt3Bg9a0
DC3hRJeWrwfSl0fuLnvDtmZZWEE+QGmeNa/FsHmG/YcNUGh1AG/+jxjkaLl+xxvd
3lKcYPERtN00ML522Lm5ZRqEevmZZSFH0H2qrYbUEB2X91jYz6EGZChCct8lz/qB
tVYKS4DvQFlU95z0/7sJNwGga2avGUwMyBYnNMv87OmSC9GLIefoGD2Li2gBRec/
cruUBBW/aHAuoSJ4lhlAIQunlg2Cz+DP8rMa65TDuPdqy35twwWReP5NIrQl6+ab
5o0DjUldEbNAJTLGIlFOMiwOw0Ce6J5jIJuplj0e1gInzi0KL3Ts5za20J93LyIP
IgSYrNDy9f+N6mUBEMFur5ZjlT8XWoxO9eUgKxuPUC65pZeFbK0QlBa0vplvLtwG
M0Bv+XqFWq1F4TJrKoFHpHQzPidBfpwFzUS+xXv4+nWnOOSS3vIHZCH6c203IGzW
5n9Kd6zOZBZB1x8kx93jNKptGSePDWmTlTqenYFjXen29V8riPXXR/TrpzeOct4e
jLyHwkHmaWsLFnxudXTj8lBGEQms2MYH+3mYILh8x6g+23uUjtG11zKJosjt1MMm
6leRcz9HrX7FnyaxMpy2tUeoF6fDY3UW2hEfJIo6EZs3RW28QBPoXQrOb/gm+erG
yDIWByomWleSKi+R1pEEYhLSxmLTTtkX97fN40ussv1oRU5RDk0JAMqbbpFqfrwq
aPEyKwQZjZInxoYO7XWMc3z+ggU9gJv8aqnBCSJlvlAsMhq00/WZ7TAk0R91XoS4
/kLCveF8E8AZkeddqJv89qwYIDKpTZNloTPMfZEmyl9IsREJEs5c9m8tGmOAzr9c
tUu97ubAwYukNsc/uQY38Pm4GrfnIRxZ2Xh2WXBw+0wzM0auYFJL0bIHcLDlsqPr
BlYlLFDi1LpPvpim0iAvAZdCxOqux/A6M/SAB22y6sPi4BP1FkypFMd0zo0XYHsS
+rbNwPZjM6JMX8xTiZyHvpXPnMUBMXFnTTRNLpOM1XLYRmupVHwfPhUXD9tF56bn
iB7qHGbvOPyOKGZQQ92OB0EjNLvNioMY8pDS+MxljuZ9BaoPC+Rytw0pObdAA5UA
y1vU0l6btjdNVr7ZSh3mR08bHWyt+xJA0YV5OWbRUX1GSK19bGseIcj7mVZHbdRT
L2pfQJlg29y2ZKspo8hSRaaHN8H9jEJiBkMzaaf2MqwQTpY/iRwVWhVD5HcWVwxx
02z5VqQ1XMmuPAKmvp3sBv5FHsOIzvMYUa++Ukn4V1JB2nOJH9eepX+21AzTcch2
+2zTLey1RF88/YWN7akzcPK7f0YRvCJms4udak9gFEvbBQ4Razr8YCJlqXpmEbTx
smlFb4EPirLacn02PpcIhDzSvAqKrquFj7Tm+k7yFBdNdw8yqh6tp3LFaF0wJt59
tZGd6I63LAAcySL2iro5VAxKK16w+a1Vh5obi5BI/n5Mve5zDlQecWKvEpj/j+/o
SdQA1ooPP9kn2n2l7Yo3v+6E1f7cNQTqsiYCeRyS/T1BcqmN8+7toBnRQMXl5Bdt
XOSy7i9HQCzzM7M24LV1a3gsU2i5j0PgNmVmdISGBUvAn7wkHO8Li04fSGcqmKSe
tGZKH89d2P39vHtRq8wfg5vur5NiKhfpXZr4+EBKQxE5y99tWuB4C0u67NhCP370
2Sv/zwDqJe+0owGrF4hormykrmrzgxt1kzVZ+5lQOz2rpx+16ISVvrQ6m1VVMAKh
+ZkuPXcEHkd2A9/HOkH9+uaCaZ9d7ZmtrlVFBG2JPdWWUnfS54WW8ljc+dUdZbUg
m1t2FboFOmHtiVISfbrgNUSFMBiKVbAxbxVHof/SUVjid77Kt0l+QFez/nT3cdYb
V16nOSu7jWCg0mnXAFFlta3T7/ba+E1yDwQl/tduVdKZUkKoNVbZh64uMPDlcRSc
YqBHs4JCjzWuaOQGjqqq+xTXQxUKK2h95MR8m9BRZnsAJ4oHRMRZsXvZpWG58uRM
771dJWqDaPSnZ5Jqys0xlzkzawQ/W7CtWrt6JGfmlAAK/52/tgyipkT9JOUdKf+p
D58a9DjSH5Hv75jUX1AmykkHQatB97eX/Ef74gNYSp6TmSwuUF98nK8pMHt0aSzm
RAA822Oqe0v7Rhg42QdrBnTG0MVHhHd8LTv8Tlit9zaEOABHCv9nih3RL9oRRizE
fOVcqomliGmln/kpE7kiTL81ZLu0itD1GncwbgJeQQLdEZbso2vKH5h+TrO2cC26
ER5eB+NUWi85BiDbSzxLYpcOi25tL4j93XSOJIF9Y7gpfqDH+lPgQQqLPiCURw1N
xuCk1ii6HGoVtnVr6DqwYnNb8VKr27OvNehiMAZd7LMdABZFqfXdlSpAZ2OpLuzW
zE2rCQbua0z/vjuIT3VzkdLk1wc/G7I22nIFUzHJkYYsLrTER2lPcANz3yPPmJ2s
Tr+p11Oazc56R9q3KZ6TZzMT0+sPeiAaVQf0OY+58FUuIhi2jxUIbLwai/icDH00
nMr6tpX00ZuUbSB9XM1HXhc932qAM3LPzqmquulekLdF5pM1YF/kkuU4mCN0wtFp
CGdmL1dnKvi6yaUo5S8/U6NGSIXCcddAo4SuueOp36YU2O2e34BZig9Yq4/qTNsX
xDKJlGRShod/omWRvkRC608jI5miwO1pQe+0PwtDjC/tekuJbIJrqHZZC38ThlYJ
rWjOcYE74TN/A7qD2gu+GRsRtL1UXGJMpQBcjQK3CLtnUKu73af7IwqIEZEch15A
rCzHWK2dqoZsZ9eVQ8po8brPTTKsseB8QaaJofjGcQ0rO6k4akfXLwFqj7elmPbx
d3OZ6QeDuhBv3mRSsJiNaesRLArNJQ7SLcPVEwB8B9ztgQWClHxK940zSIU42Fpr
GiQSqQW80Bdhmnq8PlZNddADw59JttcmjK2vRWIWdbDHViF76Urs0aw88Qd7UcRM
SpFfcDNkNdlmr16TagSONIVXk/ORP2xrixIDu2XfwkcYBxVtc2sbw4t5bBJmNhn4
JejGRAuFSndZXcuFCepSS1yYkBI6Qo0WR5Fz0o1+1N/6w0CyO4WffhOFUnGOs3ZE
zNtfNesBT/l8dmsAA4lKuDlxA8j6lVBsBorpX2InfN3qMCeXxS5e9lFmaFefLBu6
rPKUoJw+LZsFIfGRgRQHppImJVrahrv46zh/lZC3k/+feRRDF/eGf03VOrkz+Q1A
bRRR7fvxE87TKtH6tpv/W6fqC6LukRHmWtt9eEbWpoQZW1T7ZpWwiIWoiSBj8w/k
JBJZLn2oEPKQralCnckSR1lrnMSIvZ01E4v/ExjZ97c2IBk1U5q8aBRN2nytZ3Py
yAMTOY23/IvfVbRXvklWLHmimmx3aAcvk54ommy3ndK6QbzZBv5An/R+f/MNwlGr
KwdXHxSIHEVSNpHfWgSL7GahGc5a5IdEreydatD4gdpkBI/WDJqKLxRvlEGfDNob
NNZOuB3laQCdMtY3WEQf8RRnp0ZM5hugYOQ0Fu2VLVWYF8CJoWEaULyDvPdCLDhR
R1VV8+3NqsVoa0vPH+AFJH1dUqmsxk8ZpD/Dm5p7oujLYBiP2tmPndDpkMKDu8O2
MpK4SyFdzRRIs+vqaGfFnJrpYMRYBBQ7aIFfWsPWC7km0EhPNsiV6xcP7lmD86wG
88lTRvskkAhS9SElOqPg81vElhRmJjIpKtqNqyFO1l6XfYgCY4P1cfDx8jwSikEv
AJf9/PYfmn37w7DXOZ5U5GPmKKwAcWGoMs/Llq95SMzWtgOXqjzLrrzpGYWrF2Mw
+FRFKggY5e50XBCMR2zUjXTMV1Wz5lzqXa2ixxEw8HML6UZx6AR5z6KPNm16GI7R
Lg0Ls9KrgAmApBa1s7lk7vXS1VHqGHn7Gim0SlZv1fo8afltrCRCau4xHoas7EDA
O65YPKdvOh1uPkz5n20n6b4qNvHPOJVni26xWf1CqXVXmQkjiynmx/YyY6jW/xMx
of7bgXoSssVPu4HTOoQRja5cO82DwQdvDq067C+Mmca8+kzQ/2oyoswJTtHySBww
zq/G48nqwirj3GqsENwxxyTNpB3b8+nn1t6Tu2XVNGJLudkXDRfdjxmCugT0JAnu
VWljclilSu2uD8hNodVlyN+47RrZ1dxbVMM04mccbsGNH8l8BWmkpc1KTp5Y9QEl
m7vK0LLwin45Et0HV4JMOIiAfl42DeZpQe+XRurwtFUW++oi3toduaT9eKp9S68O
LJFrAp40JB0mD9G640640Gra7mM2ozG4f4AILrWsEjsD65Mo+GgiLS6ozVU3UTXr
0ot/lad6/9+zisXPlC4pVfNSnfWIYxGl6mTfHYwF8m4/jHz+T2FH7AEqtre+ZhzS
hXQLJfhB9l220OBZV4fErYvo4q7uapHhVbuUMHS7fdENeg8iKuf2e4sbxsqDen/S
vdxXtn7+BG9Kfr2ewbUh4UmjcQd4vVnH7Zmu888Jjxc39TsMHf6NCUDm6mGsGeAx
h9JtnxjI2xTWIOKUZy9sdPTqE2pdRH3YedZXVw54lP9SIA5xLcNiATUKxMnn+V/+
zsBBNVYJ4DR1HBsv3FqNh+r2976lTufuZH1wiscAelPGOcoMHDtzzF/uQnoGhl7D
qckebQy6mqk6wHDsw4dvIdsax7gLRwJQPZlrbzY8lTzTbak5cjpFgLG24pDu+qZu
aUVr1XEJd0YYxCxDeJG+dyg8XtPgZHg9gmwEvF3R9a7sdl13uvhfF1HuZOlSCHer
6RlEmEc5VoL4ZpwnElCVRJj71RL4ROKJxWPn3Z0+lr4UthHbPlDiFtuHLFYV+lm3
7etCyiLm50EbhZdedckR8QiH6/3QuV3VSE5v9VUIBrefiVr+AwMAxrQhnjpnf204
e13MIlotsrpFkFsS6DNIpW7KyQLSeO2ZSDZvn2bXrFy1r0n/Sf6+v0pOVaq0gBwn
i09801Ymyp7a1wlWk10L0OhsKjZQeDoVndxyRz9n8QQ6P3XIdRmCPIbTYyZhhu5y
6E3TxDosOi6WoPBxRg80nglM1r/b0imrL3OKjb3pP6FwkNPeGdwmsVs5yqQzfSY8
C9CTUXBwbUv46V2couQp+ewRcs4zcskj44TqNJqr8x+h5ZDl02yMRS+jk3Kyzy56
8v9aK4FUjJpN/JzSgXLT7x64pFjEL8CKQ7B+JR+rXtsmfwCPgMFelU8FQxj5mNR6
wpG7T8dcZqcXPrKR/6DuNvt6WYTVcECUuigIuwbDcGsAuSnk3ZU8C9TNYGv0WHsi
DFyeawuK7wrvB46XHEpx/odaGjzPx2qLxirU5LcoXSUrFqvSClvMrHkb88C8nWMP
4bCQZQyNCKOqvSupfdIAlhRbYyA4YgtVCX7lIZ+ZNgQA1Vxo4f5Q5sImdEba2u48
M8DBYmnkDqdjKaNId1ZFiE29TywBS+sjb1cK+mDUI5gNJfpyTyhQPivMDRItJDtv
ctjLaVCHwVF2KRDmYG+8P7J2ZLB8mPrnOs+t+9byZnR9nC4Do6mFrMLciAGReruQ
3WSUO2C9fCS9YwW2wm3TgQ5jTPXi/8k3WrEXSZTxNxZcbA8GDKWlahpC6qYgobgF
RJ5chkbFA2TTuNuLxhMsaE76fkfATS+rYb+sm9u5cZibxtVw+LgVFhJcSyxYCSto
RLUms9YGNTnDLNiV5S1kvP03y2WdxO/6PqnswICxoUJlDMW5j7XJtMNL0ahFN2cI
Emz88FWX8UElwGT3a7lUd0wUkqycBBzZwnXJa0jRYz1lnSYkEWF+kXh28yY2X9rQ
RZ0oYtFifrrUm8CUpK20rfZK7+QUqSgLhbpFvEhd5oz/5blU7jY0TRksidfq3h2D
BHihR5+Z7RBzVRTZnf+0k/J+5Lq08Gl4SpKHCchrLrYxGccJgavIEntLuREJi2ix
OKVLdmlbQ2IPKbYdM8X9c1Ia4xqBeLpjH6yIXnFp8kukP73GvOo77nEaRHkZrziA
CoZy+v9uvbAloShdTW0R9BFHH2U8PVsbss/ItkgMwAgRMZo//dUfFfrWax70AJJq
IPLV7RKjdE/ErwCk+/4Co4JnhFHgn2I0t4bIELQ1f+6KIMu6/fV8eFfkToyYHb4b
eEawdMexsFcv4Y9qDXX5MXAO+Ztl8akQU6hOzsnXWjykyTxgHRiwkmHuwJg2JAuC
FIt+n91xo/pbuBYTWh2hcb7dgCwyBy64GidSf1k+arbWL5FHjg+OjcoQHhP5nK5t
evd9z7BDVwOeR8UbcLaiddy17HAPQF4+CcspTGo2DWp7dEFrvxsvWSfJf06lyFW+
PaBjypqI2RhOQK51pga4SLdVVwTSdw6XuxzbuWMabkFelNg8qkO79gDQLFQWAYcz
UREWen0OAd17lk9WjQ6X5cCGQM7VlkE6ujxQyfCxWLLvf+REXfPGLBEKor+84+xP
FfvpsBZ8xsjpppAmIBRoWpZnihx4KaC9fpTeOtRo5bHycLfF/ED8rw2P0O46mNcH
abeqYiLbs0LxRvkAP/ZuRkHYjdFQjoAA64rExtXEHFLPbi4XkqoFtk2f48+d/Uhd
yyk9bUJVPbsGLA21zLQJvukjzK16Kg+X+/2JSMMNhAB/xFnuYt/bS0thir5haYJg
xkcWcQXL/ic/D+Cp0Ith9xxhynT8ku0lb7TUOAQyItSiwQXFMVWlbgcLeUTa7XuQ
uk/nITLP48QmrijBrHdT+hVJrcW7uun6yVHioGI/bC81+Dn9NBCjO4ZeYEe8Zb2A
0puRq127wi9D1YCR+iTSgQl59zg+Oyf/W1h8icwbTFBDV5V18kBwfsVP/SKGlkLm
Cq2gH+NNGuliMTRI4TV+tNmMbWf8LPecjtUGQGOXg9SsCMH/N1Qv//ck7yvnWeZ5
uRBMC91f7nGCLQlVcx9HhPgFrtRH7ipy1pQTiTRKutbqQeLQ3rb7+2zg3Pqu1eOa
bkTr153emB4YMCdxqc/+Tbcr+vnfmfsXcX5121gIZin+12YkQPVTXYeDfB5lHvk7
VztYVBLQu//TAEvGaKJNo0RpCwMTGhwh4hrI0wcU/vkU/K5L773ZfSUigbx/W13E
FDoGogrCUceqqGx7H4PNu+AHwbzmVMQwpqy4zrRipmwJRLRGs6VpTli3ft08uK+/
EY+SRcmfd6n8zuehNVME0Q==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
THEsHTA2k/I+mk4PxQ33vlLtRqjGurexdjGmLkg5ee8f7JTnqKtE9Lc7zR6IdQPX
7CMvGhBxsCciJKb+4qj+T7KBwL+bt0tRPP1tjHnbzhohR1Xg8db9/S+FrLD7r9Jt
gMd1vorzN5o5YP99tn9omQLFr06k5ZvMYyg9yRBht1RuzPU23i0mTlsClX7gsir0
4LsJBnrDVyqlq7X9SShZcW3iIIEmnCWlA0jTeXg2AweBGbRzXi+c8N9vo9TkB9tl
luylCDqYNNl4XQWQHPNJ/4K+QOQ3bCEc+OZ8vkj9rCdaYNZ9R1crNsmmRRfg7014
7RQwbsEumVYpEcDZp8+tew==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 544 )
`pragma protect data_block
QB8RhQVzGF3ZgP7wkFCQFMWrFJ2d/LKEDII/8dzshYx2N+5IqjcEP3HFbx1Fu3YR
EDtl270Cx2nQDXo1IW3XHgwV7nWvTit28AVgjXmgvSQ4RnuuHE8AoEwZBTAHYZBM
SCheKnSwg/zsyPFLCCk/11o69LvBrnATptpS5FvoLYioSEe4blrXjQd8y2ih9iMo
+irihGtnYwssJnUBJdNRc87hZRd3SARfC9OMeEtCjX0gO9Jz/KCm0ecpUtcdmB5P
YleJax4v/ybKn463g+ylLiCegsKzRZDNNNcA4KYKCzV2NHyQEn58gkVB1263E7Yt
Xw9bkvOoyXZnO/vvYlyswXGmeksjNowYh/wsh8FSkweywS0qFAm1Hm9raEj0FQKG
s1PN/M3YBPXCE5UXV0B3cx9aFRQavAMjq07ivnTzO7M797izk6JOzNX4Ja0i//JP
74c6mTeJ066+eBGft5JM2nJSc0vqhUVbeQBvUGszjuziyb6FTrDyiI4XWcm9oPT/
e7V+pxCpga9ZFTBMKcs5MeP2HczEJRz7gQOe+6TpLHrlj9wLAZYlCH2Wobm4+lXg
sxUNV8W0jzMoOvS5BwhZNHWgqLX8oyYOTsI0UtLNs43vEOiqoQuQY+TupdsK8RsR
61dpAjeO/KxQK0Cg4DIq5TsQBYXhU7Ep1VZKcDaV3FPXOhDOXwieAWekiU4Mqrz+
Iy/zBFIZ5+fs94t2ttCONQ==
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ED/ajCfp6sVsk2y3T3jBHiFZSSg2/zTPgNy6AVF7q5v2Jf4k8LXiH2PWHiVe/HA1
TMJJUiiIYG+DMSJNNlpivz+uXxVle9+bJfAUEzSie0mP4YeS7kcFz3ViHABc59WU
vCZYhczHmlkdLgvy/x0JcUwurPQHa7f7KvfLdKzXGcbaPBg8CTdn1dlLcYPzywxN
taAOG0KYPWgJ3UmV1XeZtfIedMEj0ShjSWViLEx0MZ10f+In4tcCgUtXCj6QnJII
bOT42tsv/++WuBA8QsaVH2Sw6czyPdXvENIsrci3XE4atfz3aib5wsgBzTBX3Oyy
gp/ZbO4GmRXF92wNMoqXjQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 704 )
`pragma protect data_block
rFvcsFfrusXuTpi6OhQcNDedo+8W6hByxgLsAkANzZM/k8xU3vWO0BXalZYEzy1I
7IThBUOjod8QtOg1x/0UCnW4bLVbzl26NM2LxpmtiDXa7BuidbHxm0JieFPhBBJK
nz06d92GMssHpuDS7EedNKcjUHW9l1Jx87kP4jd4B5Z7SVMqzFRjdvgnGPuM6Yty
Jt3fA3QGFPfyrBjq3J/txrBd9S3aMjbQprpUr0Gsz7fceJlS+H8QZS/rm8cG80Nl
b6FLunuotPsEfEK/+2Cz7O9xAbp5wdB3c2seFAxlWHBfR/dBw7ACANdktiOaZHG3
IVQjd0+DZmADPVFc0EgRWt5nMSNjwZkszXRRZUBk0MTk2C+UddZoSvvZ/caO3gIf
EOBI7lTc8DfhgfcHKg9zimwqbIcEZQZ06IQFewbUANqiAn4QMH4iKMsa+HLqOG44
JQqTRG4ZPYk1+YJxWzq8qHc5ToL7BdsDuYJglLehX+O7cvWNcEN7rTI7iCF2vMmE
y/8FXa9+opGGDMKUmaHYWK3QfDpoJtp7JrOU0jVJsDvoLTHMn6lI1U1H+j5OtGAg
stB+rarMlo+KIqUXCvHW/I+AjhrBQoBGP/A7jdlB1P5WjUMGd602lc9ICbaID0HK
6GdzC9YUFLBRHBSNTeJZVrkfDEAT1DaZyTmnWXJWPJPgbUq502SHLyYA+9laWUI9
KVbY1gDSvwIuypr283OaFX0o3pXoUFW+N3/ww84jQ7Vuur+5WKaf0It21LONtrZ6
oXRomSa43CdBlJi1CNghNgbFUH+xJ7efxCp/ps8AdTM9PePr1zHBwJCwT0gOARzk
Uj560hqGhDD8T93lII0irleEoK2Q2VhlH61t02S8mFCIz9LCrLT2v5jMLrVsMcWj
MFVcYEITDPgCUaMKxmvEJdpVa22upy0oNRfw+Hegoyw=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dQHi9qQmbysY48Hol0GfLKWDJJem1ELtt39JWSVl4MV0/v5ATmvb+r7YK9I42eY4
HOnI0bEEtlhjxiURDBNoctF0atsPLxNSYq6BOlovCAYriwWgE2YtQmUcblAiuuo/
jAutzIS3y8OThLxP3xajcWc0VoguUsBEfsHhmSRupK4Eq9j+TNamgYGX2kG2Kz+y
3OeO2a/SfaMi6BTe38Q73Syif2NzCC0FUXESvDgWWd0BgrOHEuKANbQx6buerGTJ
PzxuccWE6p2WpKWhT2iwzmH+osKU1pcg+L4YuShw7ZG5oI43kT0PD/8W/IEc2ZIn
XzRaO55EIkyz2cbQx4In1g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7200 )
`pragma protect data_block
sUm9JvrJLJRSA55UMl0j5Q+Ojj7S6QU/VtjzIC1Onerfw25fU6DqSwgfOVt4lo65
p5C2M0nj8aqiss0ffQBfXE0TDnqzxSflVBROEpFI2uweHCm5IQxnypDKEQ2lmCJ+
8qE21irtmP0rpx1DGBOPZryHfpv5UDfS3BAMusvoJdyqlinrKX8dcaqGz85S86Cz
APtSDHX3E+LavNd6tloFcHNCRT49CjjOfVtJZqFxlfd/hQK6bQsV6d05A1rxOrbk
cAiUwkjkkhLS181hLWN43VZ1BRySBs6Fhv/JBCLM+pn3vK24E3cZA3NKK+mmyJ+h
aeIj8LesIRnvfMC6r7/XkXCD09w1CWdjFDl/hLWuTHm+P5YE4Y8CfcIL6ELCup8d
iF6rde2JAdHEWck2ujaMST6hHGoViBI4lBGFG01a2yj4zFqwtKukbNefRLf3V3V0
Yq2kcd8+9duQkR372vGNyzoAJAO7MM73Gd0hHLDPVXlFyeblsFOi2sMq9AqqTMkW
OtVFZNg2zHN8My/HfR+TUYkcodXRsk4MWxEGz4i/Oi/3vhI3JnRrMdTM3nK9CPWx
KLy2c56L5IMkqyXFeXisGITtv0wtDBCnjDZ/gyqYf845ttBaEygRjUKglaiJD4/f
L3tKM8ekRaYqQUJpdvKTrOwWcZRTIi8CUUvIJ+dJm3n7NAW3dXzq3L1yulsLzbwG
5dZSCBrIcP0qVVWuIosbZiL6cdgZzZipVUOoolB1Bc5NKVz+B6RZhqW1e59SRckY
o3dePWiu1bzShDD+dc8MHrn0sAPCkV7w/r+46Y/bZK4+C376cNLK1/j7ueJFfJxz
A3IZD6nYsyyZphnoGQNlSSPFT2B8wMHTHcv575ffIaNel4jZvyoSLIVrZQwmDeaH
8hLRp1yCb8BSJVQ47rqyz4NrBUzO9sp3tNx0tLUSZ0uPWEF/G33GifYDIDyNbV6S
T8tMcLPED/sxMT6lcz7LvYkd2fR2plsU3gqVzTglJqPxlEa0zg5vYwalSOkFzf5x
npxiUuKJJCe3Ghn2/zh4ZmOEcx6lYRdz1Wr9YKbFTRTcnfu0R2OmWYvy5+N0E4A4
+oG+L0Dvxb3brcK2Ydg6BYcRGr6ODWt07SjOf4RumPVXWs8OVosL/mZVLFfT/PBs
2yfq7UbXEhU0ToSyuErDHdUHkZueILPVP0KnellZOMCyAMsABrEzXaZCBRX+vOHV
yxwfeBWQNctusrKjaNVjKExtMae47mpXlet0JDD9bdyqpcau0JckgeVGXme4wNiz
eMnBRY24qcqgupsN+b6ef8iDS+xilSOzNIhYsHVy9U/A6K4ck6FzLuNKwuzFhhJ5
e2b5OBP7rTGI2N/3LEY0RlVClnSlJ8FRkzT1BIuQnLBBoTHwZHZaWYRsqhMw6Ed3
xGwPKVY4MuKAccdoW5Bu9yuWzIdp/HX5yQqG9UQZKob8XEpYns8qYbBAltG5616p
1coaT3/y+GU/oRQeeAs6YkLpOGKn5DUMRjfxM9jfC7/VhVXNp3xqP5BizuRQ+liU
KI9bWcdUZWqOtN22A64DlgqqMP25klxike2S6JJsGT84zQyFMcupMdcyMZRO2d28
EJHT5DcaTeICR73NsgVa4d5FlXWjzs2sr5fohzY0cub52CeHt7GM7l4+fG8y1hw5
zuEGHe3U+eU03KZ2dK4NVq0s2Svvjsb9TPSIiKqvRKhlMWgOqK3Km0RmmI2s4rWo
PTTjKyKkkj/fUsC032vAriRcnyf2ZA5JhXnClSW1kxVhdsX2GBKenYlifyBje8DH
yBuYpM9GrTrWr5oSAvHgFXzSIqV2LNyozzYUhPbeV6OkmY9IwH76pEgwQg8r305j
s0u5BSUOepLpL3NfB6G3YQEAbkCjSYAYBTFvKDtJ9WmaWVlz/kOueU7i+PuEqRKb
pGE1g2jitI5/oZlIa76Lvipb/vJqLjhfDfoy1YUzPFIcqj8M61WdQ4thqUzLc/2M
Va/bHEUgP6dUMon2hdsLOQfUFrr/e4uVJiAqIrWjcixzG+oQ+NbBNfEGZnLjU7dt
+L/dbFRZP/wNrA3y7z0L5YIm5AbVIgYjKSohV1cyT/eYjnvEIhg9vHZRANlYns7d
Jtk0yC8atVBpM8GWkKdAiBscR6q2cUuxZ8qg8CdoIDPdHtAcn0noh+21pdjTpsFI
+20KB2oXEqdMXqyJ4lBpG9amsJEOXORhr/dR/g+DvN7aZ7bwqzd3RYoymuig48b1
qpKsn23j/57zsm3PFX9yaN4oC+nlrpX8/g86b0zfaDkAwRS61zBDUPGA3gB7Cqdu
wGrxMJ8wkl+DJQS4iuy/q/aCz7PUBse34cnnxXTZduXoIf/Kz4q0ep/kd1+gAzAz
NbYvlDtTI5E/qwX7wT0mDkdGKn/efxV14ltxFRHYNo6mm633JyenU2tAlpnq4c91
6tz7SC8HA72zQhEcL6r52slOW4ED4u36wT5bmmvVBqQ/dBYSXnHje09KF9vcttPF
AIlC6+tZJkWtwjQ1daC8k9mS7oC3AZ2NuzfKe8ob9QJw6sH1BGmLL7yoeaomX4x4
uXo3p3KNZAkGXV1k9jpRdiV66SLAELFfTXd4G7Mp74VLoiwpvQQjGVUSV5Dh8eiG
df7r7ZvvtNN0175Xid5oELgECfFLKDVRSAyqYmwdvgb2DJqbVcSCcMk6AwRtFuf3
OEa4uBG2oj+eTLC2YXhznp/ljTGerVG2pPqdJo5QPJS/cFbS5chmRDOM7CTWd3GH
/mBWuY5ZBkitDOMT4xxi9txQzJGkBoVjLkfjpDfHP4+o7S/KDcMhEOU45u962eDg
90IBInZIlHdYaqYgDQKw0/BwezXnUEmnF3sVw0g1rkW9A95OM3adnDR/l+4cVPZ6
ey5nRivXEjjkrZT6lXM5yYmsyjcTnek3ReI/csoezVhdjvTq/NVgpMU2npCt9DRc
0CIAVs2oqvQNCzCe874ol6nQ612KJZg8FzSo6hlG/kKLxOAG73JJniJpuzR4PSNs
op+lBlfZqpPzWntB9+ztBcUGV0xcnDgBU4auzNFPavAr8b4UZ7OMYhHtF8M97X6R
wfHAO7puRywfpBEjI9IME/Aqq7i6DVN5rQl0hHP2iklLV2YqPxLrcwHMpzqO9WtT
8859sM24fQrKHNAyQW7Qt9V0T1RVc0ZIH68jzqZC/GOP8+2clon/DN3ReS/lLKB8
bcWR//T1OzQ3ANj3syE6jYBaprOchSPB+PIM6GDlTae5mXJhKdR6ku2HSQA77+DZ
wvQiYJYCqW8OyyxG2q9BI6C/Neg4n8TaA7Np2TQwOfqDS9H5+Idd0rP28AMnjrWu
9i+wdLrjJjwxb1Me6HT6hJeaCdS2K9XTeuJQ77YTnVgAONYs+mZPitoGpHOQeOhW
Rm1nXSXAgjD2trrtxCbScJe4IQceYgjwTKnaEt7I08QliWf9WB8CfnY1f7UunZGG
p4YgC2/sxD7nTdDkaW0Tq6pLopyWbSHZ7iU2N7jFJqUVxcs4VFM0vYX5v1XKq0t4
BQNfNqAz4SvGt2syHf7aqkp0V9p8DrILkzmEQINeZoSlJ4sbmdCwG4iHYHvp8uOC
UNinM4lfpvPEqpCvrBVRKjhIM/752OdIql+8VPVnoGnFhqFxXqBxuc1s7uDRtpXQ
sfTQfrhPkbGjgNO0qLd4E4QSidZ4VxYcommmM9WtFLC1Afe6Xg/xLK9HomAAdYBm
K4R18mO0iLWiO0beXjZqQsiUr6G6G+K5a4ycjz7M2gq1qINW+I4/l+U4EuOo46Pn
JWC9dfFLCnUidWflW+0L/lepTqmuJ01Exqf8NJyv8jH0Am9m6Hzu1roPC0FkzI/L
8Y2lBuG0C7eCTlWa9b3FgPdS31IxvGb7tjLR1iWytLk8Poes2gBHpyksqZDO0I65
FXKb3M8e+ePIIKN9iubNVmUJvWsibJ7zQ9P1l5OswOlLJ0vn3CssdbdD0ApPJa8O
P9UiG5YU1esQ6GbK5+8V/bXTjuirSMl3hQr5kvVqrl8Aprl5JX0l9NrVDprpJd2q
ocr42YWvAXyGFr4etSBcqGaoe4YYOBRsj2HoGjw21/E2DPsbjuiQRk7fSBxDjjaj
vWHA/MLBS0IgIDV0tu9EjP7hDRZZ9QaWbTT9A2hzEkvDpfNcWnW+fn2wgg95OuG7
fd8q3eEfSPgP0Hj1SvPgs54OWhJQsvpbxhTlp+dAAJWpYVLFNMOZbEcvVQ3sZS+h
Vq6cQSNPn1FRL8fZ6DvhrGDGAE9SQVrpfZx1LAZVoI7CkhS3y4I0HaXomsF4YUVe
IHhdf0dGkgHbbD288OTVMIufninqC5CHE+4z0jyaIz02j9hl7ojaMiRz4VLH1ie7
xFGQ5wbucmsz/ZRDJ2u/LqSMA0lK5Fk+7dIxijNSe10aYAiZ0I3xzMQI/NL6Niq8
VhKt9hi+yssysQ0XExgOqQ8l4mMTWMjhARxYKJTXqHISsTkcuQoi2IZPVExLs9By
gBcuFCZELX1nriN/NDBOWw7ZyK88XaqqmwErpxIc+E0BJYJGPsllNo39XcYu1ppq
RS1nV5SJxLl+B8ewZKb7E199AEhh5F91mWKWSHtkpG2hdeb2XPrDK0gUsEfXrPFy
p5R31f5xU/SVWAM0qLGJTnrss9GdIQZHtobrvegaa5AdZIwebjTDwHmRS7Pt8RT6
/CajXIj/GL1CpFjEEW8E7bmAh5Ao5SDWMrn+Qn23hlTuh1PzbEEAuNJR4Oob1HtB
3W0+HCsp5WK3+Kl5SA97dDFBYM9prvYaHchLl98wuPf3LykSYT0HvSpSEOSEWbdy
ZAEiuqFzAkqcrfkgXCNqJR1wplYEgOR4khFheZOTetMbgT6V9HafadmY/dk5Sheo
F5ZfCshfAwP6t1B4+lCyEsHPkkWN4eQQapqfulTW7YSN7IFII8G4jc+YB+etFkAK
7IQoNBemAGU2nifCnsJ3CvVgtK6blIKHdSjG7t823PAGK5mXlTKLQV+vryNatyEb
l3x/hkkwdmBXXPnG3TM19fW6qkxmN/A+IRqipp7YoTqkR9ifQWXwZiVhTtJvEej8
vlA0UQ5RDtJ/qNTi7TOZQ0WPA5bn24eR7hkPriwWlhFi6u+xIBvGa4Sqw1Lrku18
3RV4247bSUfhA3X1zB288MgO/qVaTTA6V5CIMAQzYyByhCyYJd9ZUceXnxdXHEKb
Vkmfa19HG4np3XSUdhr0heHEjNbpvoSAEj+XDs/EZeppcevYbRjLkoMW1Rag9G0g
yLKbtKW2vH4Hde38DG21/LSmiFQni8CEeFptkETVB1XZTsmryEQbN/nuakPpxPno
D91XwaTGpW/rTbQILB0B+FO6WfGUxpTArFjiTaITcBA93+Ppcs5nxqAc6Iqyp38C
HkuRQTWIuzykzkGiWoZtTP0JQ6qfGLKwsyzYFzBDTywpKhB5PrV7loBjuBHpqMUd
CNXX4clWBSZ8KkLmD2WpwYJYCla6qE3YL95VMdKRYwO40tI03EfDHrHvw51IXb2f
FxCslJ+SqKu4iIhhEOWS8PiKdQAS06EO71h7JRlF1D7qxnrZszm6p0ZA9Sewx6AZ
IiB5GCvIo1PZdcwOqrnEC5iINeAltYGQCrPS6jw0Qi13G547A9FEVYa4tBRtuaPq
TE3jv3NCqhjpAUkBn6fngPWBUs3torV/mvbBu6GWWhOxoqAmj6vXPrquy0kAqmmX
unvg+WfeEE8/A8NF4F56bMNNBt7jj3pyM1UABVChGJ2p4W149nL/uquUuv8XHwW9
ceA5XWQ7e4TxBle/aQTiLzYQH840iMbM0/s3uHirYLPit0zULqUJRhK1bWl8B6f2
fPJfg5qKV030sYlFMQPdtVfocuo+hrRxwNYh/ttQZ5By1fUfpaiOHjUtJMcvA42l
xsfen7A7KqiIj6117/qNNcdr0c/wfz93bdDpFeDGPiyDZti0y7SIijq8JrJiXqCv
2zsdPSb3NPF67a3dKExV/yZ/SEyCn4N0a/nz6M7elQuWZCp4nFmlB4mCjApXNjpL
vASZH2BQQofafh7444r8CW/pWvn4sA8gpPGvai5qNRFQOUmlTbthFDLhURbt2rWw
KDK8pNqmqpYRXbysvScOjgkRV1M8issV4xBbwAnISatbzqMLA4G57RcrrcJrrVwT
RRJzdK0U0JykBog14deSWtxmGx8rtu5gwIUWvpgP4nCCSrCKZOIQl9W73KOk93za
pKG2JQ9toQczWI0lGVis1tpZDLilp6mPrKFFm2/tmFOA7W98gkpgdrSOss2aKNfM
4Zufn00wgS9w97viY4DhiodpwFCypK39cn8coIjcR4EriCBva3+GBXeH8gzxMQ/2
iE3fgPPBX8zo5UlQTf+LF3/sGqnNq1yAB16M7z955XWUi6+Y4AdRpbfBt7qeag4I
7ihQrxvFfY/2K1D7HztA4NKcqneKRqJT4zn/1HmlQoxK2QALVnF5e4uz6mvRuBRF
4Z6V1I4vOd1QcfWtRw3fkEkjEzpH4lCarSo7af56DAntA4Et/Cq9Bt2lE2b8brum
JoGDMU6n+XBgnXY0bKLiY0XmoWGPb+XVj06tPkZPboN6j5RbyT3aB98mmNiC36z7
ABzoJrwFDTIqS4KCTGBtgOs5d2cy5/T+7d1xiTtElJnzWKGz371XMLhsbQYDqwMk
T3zsC4oe8s+zbz+NuYrZyK1Rq9kIkIWv1U6wGa0fnAGJud0OhvwGJ7f37QgjgA5t
GRxpu8EMkjjMXdJ0uc0EYFcXHjg1Esf/pIiRypR01T6da9wUT8gO4Edcwr9el48o
ghuTdRIdb/p7zapB4OpoQQLMKyD/SLgqsNnHjKCWpOqM5Jo9DxO7i3CflUs+j4xq
SDwGUhVggD8rQDNczB/7DOkDyJaBZXVqZewSZ5/PHO5fivOa+edJD1fHrtPLAxxZ
rGPI6suTBy/nqoVVV8LWcxNdVlMV8kgOkMiSz282qrHVtCWV95acobAOjZpF6uWX
eIzsu3yCdoqwqlkMrKN3e9r034JUh/hr/GSKpWhO43UwoROZ2falyl7n4Ya4cK+y
6lcO2KC/eLASDYIcr5ymDZI8fqsRnluFALvM1fXwoWCEK3vm2siyHYozbBrLV3ou
DP4Et83e6wf7EnWg1vkb+SoR1OFgzq9cqTYs4L47j1J8UoUXFW4ALlpQ2+W7chQ7
L6/gimkW+nzRb64khXVHw9Lf4yXGzo/gr3/5sVoeAb9vPffn0N0aUjo2O/vyv3le
zgD8EuozTXZ9kbm55jFKYkYoULDkg+h5RZRzcdYTIu2uyWu/CAkQSfqP/IIyo6vR
Dg9i8akiV/IxUQc+oVAi4XUvN1GlU6s3QcXoC1AaE8pL9Rtz0EcAjqScSxGWjVHB
5ZbnCmgqyLZq4cJ2AVjq6FxUaWPK2Bv7tL9jn7YlkeUyK+ya7nKDJ8TUldKGX3GU
joV1UobfI0RLEsWMFLCNzBlJ+66Zg9sjhsLBsGPyw8Bo4IZQRgQy+5hP29OM+JE0
kKVMZ0D5+6+iXPo2DR81rO/Jwtz02Vyk5keChE/Jvu+GbXT7Jrg2TF1bzXhJrDpX
hF0QXoKp5/XWJM9Lq6K9/BJi5VqugdLOeAKJMucdDwbHEpP7EuOjA/osIWHwVzcc
rczyXoQCAB7CEtRGPpiwk5Dz0BjZ+ZGbg7tw2LsV7s1uBFug7vJKaQsDtMlJCPAM
ndSjE7Rt2/gFmmjQ7PH0tNo4wdWLttPLRFIamzqnBmd5ujSMPRCNtIchFP9itbvQ
8n7MYBZ6Q82NiueHG5giW52w/wGyycVg826bq9kudEDxDeV5yS/BudBUDs1j0Ous
ebyDjzYM4eD2ApAk0WigUF4pgmnPDCUy0Kvy9Gdonc3EvR7UrAefu2kgpTcL9Xs3
/JHMCilziKGstFIAVZAlrUWuoubyBgMAwo9Ez5Q2YE6kqV9g9Q2nQzPCLolJqML1
IPk5yYs8Kj+zPOt1taHoRafr3c7uUL9g4vGYpnnkrJmNV4r/4d7N9ptDyJrCmW9E
Ke7Dnq4YBXxAejJnAAjSv6HH4Tv+T6vb8bDEZ8cxs2uIs6/+giW18aWS8wN311Bg
f9E6eVvC82qNl7vW/Ynd7B1NIFkUt5gpdSBAM9Lahx705O4w8dJPLVFUkMkAyLUF
t7rzFB/e+rN9LpdlqLdiBnWQz1DCOhq6O/TcL6ikYvBLGBHur6Mxk11KTd8vVV1c
vm6+o0+KHA+p928PBdyqHsWuz6tlF7j/SXTXfxXM7Kdtg6Uycd+6ABg5I23Qd5RH
vFNHQSu9xEGJhc8gdStZVaW4TWBIZfaappe7SLAiLyJrWpmLRTxmcOdeYmS03jmK
JTIHMwvWWY7Pyl0pcc6CknLdK3rPbEeZQmSa/TOpClALX3kSmmibCcv82EYvKdo1
pTtm8zcWBZ4djg0tN2xZgKYaAP1WU8pVaJtWjaUnLVJVpIWUiI4DI8LNMUDIsLEp
/1D3zvd+9qTIz+qzSokxcT6f4Xoo0f6ZZxcWgBSPQPVp1jGfviLwn8H/jS/cafx2
MnWqB19nqbROIDvLTqBuU22f4nDkgyhWghx3wlcmxaCa0w02iZzzqkRyP6VE7N76
cOWOQ7UhQLny9ZAAOd+sXOrIe2th9xnSr9fb7e+mo7AXfBYSkn+Dh6/sFCJqvEEs
bzS8lZta69sOC9yB3uuxMJYPG6+4d1HuuRyYPpysopDOMoGC1eciJi2FsT4N4EnD
GkoBjByzkVc/SIJZB8d9ncRefRIHj10qR6CqS3tKwKMqWFdm9HnWAVNsJlCe5Wqj
eUFDaLap3beh0iTv8LUrNpFgehoT0iCcBIglH5vFLyxEf4/vW7GNC7EaZznz40Cz
ZDAZAQR5JkwqOFVNpfMxw4fe9mxpZaBHkstJQR0tyAc4mBpNTz55cIbUT8+8inv5
pFAjAPTTT42rqTTeCphA1nSEPeVuvCRhHeg6kBpJ0AzMTt9vui0EZdM0pHmzkYh+
CmLK1gVm6HEy21XgSJEqDiiRtFsP6S3O2Nwpsw4IAT6CuWAz8SG1S28XVB6lDxvM
hJQpqiJqQkoPHo6jp3DtvvUdxnpC4EBiNmiMm7Jp0lxe6rMwexdztk8IAJJ7hm+K
GyvNJzAfBoIzXYW0ammUY6zyhj3rbETV69Xxuh6TKyWRogjDiUv71pnpKiuT8dU1
5n4JmrkCrEamtcUBE/uSmGKb2nGnD3XWqzhjTwEB/bRt7K0WQ6xvvCHdRxTv4DXq
pvaOWHlqk86LGAvEjZpkbcRBdVACKnIq8kdzoLXW18b8Vo4yJN4oxf0Zx1/Q4Cvz
sWZurixDb7bMouTovuZxm75Mh55XHZx6Hti8FjQRqH45TGUzochzP0+uyH3EuM50
xDwjgbqyAQgpq3aKNzwd1QFsVbviSMW3o/pJP+3kUrOdfQVSE+F2FzlEkDuEaVzg
94D6jbl71hbrMVo37TFL8VBo1KAUGj7rragXRBY05TlSAMDncpOVWcxURosUWvc4
aJq0lu0zw941k8WFtBBsinGBYfocGwq42S4LYm0u0L6xG5oxRwqQZ+LH6Sh86/CP
U3KmnDBpQkomAVuhKjeMqJ52NpdD5tUCX68KrChplXrH1AOqB5GgCnae3Qwv2zVr
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
CvH5XodKSQq9YmGRE5IQW3J34dwqubvQQ1vTLIWgdeMZyRbFunFEC6KlLeFUUKdA
V8r3k/xasTTMO15ZF2xwWLC1xo88sDkfbcJWg0Qlu6dsacyKM8nXRNK4GTLv6xO6
uHTN6fX+5AeMBDgfAP3D9V0AsHm9ftrl6u5hHPoV66e0Ok3BEyfXToxo/li7sUoa
eKeZoDiSj+YZcHt+VgltqL90Hbf31tk/BeNUAUeAr6K6881tGDwIE1x/Wg3tSs51
gHrv4PdCILdpS170xsdlc5IKEHiDbvVc63dOK2/GrhJ+xKsQ9/lUSrgNzzebD9VY
ljxBLUqHEjp6r921JO9mKQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9296 )
`pragma protect data_block
pjBPNjmN8jQ9sjauugvMeKAiZsFGEr7W9ofYhqkBqN54g2f0+e0Zz2b9p4eAMSGJ
gQ8JrLwTQxv6u5LaLO2YDydayFuf7WovM/76b9F1101i4HyBiKsN0pZocw78jzki
6q1MJ3wx19FOH5VoUt0xQ8O+70h3yx65P/xx/qUQM/+HoRgNnwAAfeR4VzlCk/Ic
RDKoh+Awwb9UlSSoqb7zWRhqgQ0ghUodypRv83cM41RZbracHYex6ZGi3mplaSai
jfM8WwzFUqKb+vfgXfQ7uGcbpeAGB/DysvqTxXOqReLJlxo1llqRr1beIo5GFC6+
LT0AAUIYtnLtHhE7BpN9RucgePwW5vY+aZknrxkeMjEQZpXCOK6tL17weEciJRUC
4KyNmSraJoiuS9GwRo6VflB8vj+zoPL62o/Ij9sU9qsSvD38TbNwa499FDSGqJ9i
H07KGNExIE8yEhwZlDhncYQuDX80klwdplIPy6gSqP4q0D6wXNqsfJ0jp0tOJbVv
QuumGYg8J2Saorl6dQ3ZOsuGgYd7psnVuyN88UxB1p88VdFrwN0g2pOUfDvvDkNl
e5OUT7Ea/evOwoDs163UXiCepyVOej7YXr9Yq06U9y/uswd06gLtcn6qn+yLm1Qv
6An5xk02wBJBjsBBd87Q8fUXePu4xo1M/LkuRXrDoRU0Zmivd62LzUO895uZ7U9D
DS6R+EtUz1bpVfXlbE4TnIN/uzg1C0Z5qmcmTh4hWYpNBYo1Ulr2rBYMntIBSEUs
nAgOb1+2kj13nf54IM8Mo22EjJ5Y+bo5AVALIlhglVRtuD7IsehRVl6RZnWRAkNb
7BZ9fTDMPIaW6zWNOBw8Et4SovPoAyg4ZwOTWjAOdsjp1TACrnbRoF6E1fb8NKAi
Kes+2XFWRUxoACyQ9NtZ23OEPrDP2Xubxp0ZgGYIkQ30RswBadbYRsOkYF/n36KX
T4JDIQZmYT7+MLHqWd/caDCGBNlVoewA0H/ybC5f1lh3fc+WB3Ts22tmeKZSLiOg
DRpBI4NSC8+LX3E5YCQirv3yjnNkIUVKKFzJNoS687aRIcvuUkTMvfkHzHSyS6is
7C4SOuZHgHarESB28RT/g5oVmj1BA2YibbgmEIo4yDWLBQvzpV+6wXvPjcNj5mXy
yrb1+ZpA9K9d7N+HwkTg5CB9RNI14ajyQAOV6qeJt0Vey0xIpiSgdonfvEX6Slli
vOFoyTPjgTUkMW2CfMr72ymG8XFDmU2DaRCOSY0QQbL1sypj6gtaDHDwheWooOEr
aWbJVgRp0Wk2+A7Wc2eivQDvyAVcRlRidswpk6qhIYGM9E48ElTKT1HUbDWUK/u8
Vb66ri6G18aJ7Bi5hvfPnEy4nRzvlMmCft4yO6Yqji8mFox8LVZ3RzZJrsoq1ned
KufItBxSXHJ6i2La4s5PVKjC76XoamweR5/ydx2sq+fDby7XfMOmp82UOcX7uRsN
BxH+/1S5rBNeuGmjfpVJNMIOHJFGda6BkEECH1130MhxMGhjdSSFxqZMXblsAyvp
hJ4bDJ3Vw+aQh4fJdaU9XlDCFpN4sB/cZQa4xxvJnfoM2Sl7KA9GRarxJ2Ih1CM8
0hz1bUY6gOkUgZSbDnBzRryIj2UeSOXln4r2bHpJlJPuqaW2Xz8ZRIyaXLb5CWBW
cUom6nXqzh6Utz1Y++CadozHKaHTQlLJDMJNCj+LRG6+4S7tXx/KsOaNgbXyn47m
/Mw9Flgu0ONbX3gZs1FXUfcAmeASeou5pX1xC8vrDkMQgzKw5BHaGkNBDhV9+m0v
CG1xe5NX6EjRea6QDpmUf+dLSzphSUdN6hcquEezuugxo1WYi3iqtNA84kiWQrWS
9cragPfGWd78ww/MhEnBasxLuVfpKhpZ/7Blb82u0C3GFP5KD//PkUt49LzPZOJS
pW35L9F1CkqPRYrHNSFufTykGqHhpHWjdXhyKXyCEMgHJIs9F4DLXMx7Bm6pZU6c
Lf4Lsi58zcqLwYl8weGwwVVI3p7JdbnRvUC+1CCkuaDO/raCNfuFvHsIMwa2cpIQ
/+xYAvlv4EF9h+IspiM24+V4/SY5/vFkjxf4tCev9Y8TQMrzBAcmuSX1wUV/lM6H
F48mUhfuThI1NESbG8byLZ3nYPL1ZeuAXF7M+GXbLmJ8pLTOIHA9N2voxRbmgevi
izRP7CxByxazPDTcp0hLiThKnxrZo4CYFn0RFjl9CvaompKlnvBHg1/VKJ3iaoYg
CLf6Bz7SkqiHNx+iK+uQv6jm2Rq0IQz98dFDUXM28ABIQ3xPlDROfRFlPb5nnm+L
yEte6qlE36WANO6jEH4oIrFr/5tIuApfqgNhYLYR6gjYiqXw+kiQzMAFe432r5rg
F7fKZg3Op/JSLwnBTkUF9pPol8OXOuyEqBaIOwPeXGzmPr87oYR8DEozcxephclr
kRrtoJ5UA4siF1Mqi8rwG9Jgrtl/E6qF3FAahvECKl2xSkFbF3KsyxQP0vCtzUr0
Hd7vLscg4b4SNb3kHvDJiPiumFw6WHiqa5rLT47CbkyZQmV1IZMg5doXSO6HK7xg
HZnYx+tl+RHxuDl9hbkQ6wCE7jVg+mGYzVCgEopaNhYB9/VD9ZOwHYJd3mmm6V4D
J6oymlXzwBcCAI6mO2G7RRa38koK91/7skR2MBA+LsQKTYmfUki+oXyDOOsPGD7D
I2pGHHXIPduC8XYc0Q/zoyAnUgmDp3+V+4XnhpE5P/5VvAmkc7DwimM56mCg7rQO
sjGQGCmsx7TI7JWX2uVRO0h5O/7LTeYx6zYbWTcX8zFuwTEcXoixQFS97XnxMksR
WBNHSglLFHORFvAZf9KOtiNcxuI5kQkwT/cu61hrMqVXSs7715bYYXVWzo7v5ny0
yldWOB4AiJ6xH+ajkRiuEDxxW7+Jrr4S0dYd0bsMdF9S942D/ZhimqMiWuY6GX55
XQO1eobCtlGyq7aBelSYJ7j1Bcv9+GBJYb2W7HwomEJyU043do8zSaIVtHpSQbbe
tMRchF86yZy/un6LAx7t23vVxAe8PcTTn+hWY5umYNeaw5bcDC7WhbqrCiAaxY1t
2bij8fUs0dSMpkzs2+BUDez3O2flnDSPic9q5WyQDLa0qz3IbMlmimHcEn+iYkWU
roQ4grFp+P0HejjAK1JudacWkZXndODTHRlKnlkeJ4DJdyz+2FqE7UDKum2I0gzq
6BUuxxoT8bf/5b8cRz8zM57/ayE6zIl64EvUk671XqzzcVJTX1CuYEdUApLn4tEi
McGsCn2DBLzpMw5QFYbvOd9OUOvTnJMH2dXuMSADv2xb1DqCLYxprAQdNZtBfswS
Y/D76UhpnkSFwtUOnyf0QYWpyhrc0BvsmGJ8h4jRRd6PKGOCeQW+j6/Phr329Ok7
Hp9ICLduQ6tvGx9GLMPBwUKbkfw9Dz1lvOI1Ven5gUJdlbLkaPypN+T68eOHVAGj
KTtVWiXX0Fu+yzODQ8CqPXOHjtBhPIAZWeILjgTOmxL5BPAGGjV8z2/C0SNQyE8s
AsKXEIlp6T02NxjsjkK5L85OwgXdZyCKkBxQvFWCKJbQ6uR6FxnT+45QC63omSMF
3uC2EbscXAmGzERCV/ABk5mUO++d80FJOYTq3aUz9TwWvSJURvqNvkzxngWKO4mh
aChWZi6G3jPZnuGm/A0UZmmeZtwkKAdLlpegCbmZAzOnNvfhnPzL4EhRuOoxa98r
tGTf9mKMUZkQEvyD0UNk12TyThkqM9gzMlOOCWgN5vuNbqIxjCmpmuZA9nwzwkEg
FTM/9R8V45wUlVWrde9MEkKyvCT2tzqz14/J4I/XmTib913aje3dLL3hKrlNkn86
6kjcUhdbk1P78x8ZDovc7de3C2ScpgNbIXbhopOBcSLPlJ8CvJXz6Zu4CzGEbd1i
Chla7+CUNH3teyiAprPpz6DLQw3QTJHvTLK8ZO9PTmF6JYmZGPU5ZXQFSa7+pP94
pJCcnrLmMjfVQhxN5g47yc6o5CIfiiVDycXnA4nZII56JjINk37Gi7jesN9Yt1ns
hWV67Uh9Auf640otxSCCRv1HM+2AHjNmS2ulF4zqJxp16bsXkJt0WmOX4X0/mWwU
Kwe/PkjwXm/EbKgrHIezyc1iHO2qBLHZivC++qoykjQ9pt2goJEo0jMcNUF86/7O
W2pznMKthS0gJ1m6qdZiT0zXpGWZ4NZOxBAdKoi5FrbjSVipxo9ozM8+rFgHGu/g
9WyYtixwPDbNpoUjPGI5oGyXNULKjfgs9jzU7BEA8TrYmk1kAjvYmNcAWPRRVZX5
oQqmfhVL1adHUzpIlhqQXICPzK708gkfU8dDNZzz1tIcG6JE/eznPWSMiit0ah+S
Af/OiSmK/UJcLWMa8VMSDYPwtn8RO3/iVzHMYH1h/5yDl+7SULWeP0l7O5rK75oH
rMTbK63XjwEBd+bhmo+aW8HrLkwJWQ4pran9TOfQOyfaF9uV8gi22qpdltw1tO7W
+Qh46cEw/C9Gg3/uMryUzZED/epe960iZFk1JOb+qDLPasLe0y832ZjJxigG+EZ5
aA/KRXywQfFUNq+DJWpJA2OE1zEHOg0s7wcTinbGrTVelUfcyKGecE8lTxmLvSak
uRVlCCcrvW7JEgCvutIs5NXM+M29wSl5R0eOZJu/ZVytlmfYNmB+v8AKZUJe8yHD
cewV2p8DSGZ6A322zRokebA0C4Mautr1gBqLiR8lIc3BSBhLO8rtDU0/BfCM1wc2
NOuDYjgXc9xlilwwRk+kkLmeW40nxwhtr+UZRHWIfrqOYS/RjJWrEB7Qzvjtly2+
Chm8lThPgl4NmhDUU7FQzkgHYbMngZwfXrL7nFJknlBdRy8Kv0T6MXtmo1t8e36s
SWAj23IA86TTMrLwsVCqj5W69DAq867/XQn+T09/XH6m9VyuojN374PHIs5G5pd8
604oE7WhNOGcRQK1gmzeSwYgBUQb6Hk+QWah+dSxKOJDnfKpV661Hq7v8SM2RIYG
F6rjsKe7MB+XBhYv7eriNzwXQSfYCmmMMVaI/b2BHlWjMOgQA3JUv46euINJZ3O6
acDWqjbYkRHPdBrcDlswfr4ZKv25I7UA5YgQuebg2KJG4Teu+6FPCYaY1Y3GJotg
6FTnaQZVpl2GQXLVUNwmkOy6aTmSBf8xdJfTs/me9foyLq9ir4dHRTv60ilQhuTz
Ht7aIVOy2UBFNZuR/DanNnMONlaLf40Mjb81HdpnvVlNrgUgJTcbgPfmBPl1RWlk
1Gjj0GxWQocnAdov8h6rwhZOfZ2uMNH6EiYrErJLPCaGISYdtQeYCwr8khezzm4j
mOvb8IfKRTipdFfXLAN6tLOfWeNKOzgqIdgHBST2FHASTTpXSAwnV2G/I7qsd2/m
5cfnpCQWTOJxf8iisqY/8JnHi48g0yGMH4ZmRdRBA1oSJQo/H0Cuz1Hf5XKzqcyE
y5bnwkfsU4CposKEkRkPYVP7dD4KK7v0mmuBJArv/f2/zuaHm1BQPb3UjHdiJp2V
nXB614RcD+diGUveTN9ZBEdT93F1cpAOkK9L83zc030cmVIDVI/cd2g2SZ2Lsw5w
Nuu/gEj3vl6YUrs7s0q/WC8w4+B+3t8RwxY8fPYwaKMUeUmzvt/Y8eZjwPfOM2Jg
fkh/SFUp0QGyvj6o4OdNZsmOpaPRbggilGrQ7QkKDpOO8iyVYuf3nlEdqLWxu0Rk
krFi148mLxUseyJ9eFkHzQv7LpCEHcQBV6GKvn5KVbDbhnzQgoeDjXqIJxJDFXe2
fJJezJQmUHvekbY/oDaN2j+Mp7LeVE5DGUb+bGaDIbdGUUvUXZNofAgR7fPVOUrQ
JxMonrFXPFl5lLX/ZaGf8DJh6B7d4KHlEKhs8VqvQY7idVtubRz3seblV+pFL9Cd
b8/PyTfT6ZxwRsSQGvapLUZYBlCix4mFdrwQpV9+CYeFfdtoDZnE54MXP5fRI15+
7ccNVKUKGMZP6rtfmtjNLF8kdgrKVYkuGakhfPCLujw4a34miDzyDKlahhgXMt1L
LXv0YExOsyAXWWM3o1jUHSiisJo1i06D270iitObNNhbh6cPC33F2+awC6RzblZ4
POlBYTQogJ8i+mHXWMEKzGwYKYJsw5rOuci0oPBt0ri3f7paZZxTps+Wkp/ZRJnJ
unNlONef26j7c8vQKLhLNzEykvvKBR2/pRZ+VHdq4IVxB9VOyBczAyG84nMZm7ED
KuHZ+1FjwSb4GasUpS89xnES33ah8h+QusEqebV1p0LpMeylv9gz1BxA3tg2b/z4
dJaojBeZ5Xa6Grl+5mVVaHoFKNI+5EM+HLfgqqXWf2hbMBAJblsGRqQCT2vznWti
JfpFjEuFtFLWasMK2Y9UqmBMOg/hAy4ysEXltmdK+UB9gJn2C43+V+hz/1fuZfXi
CsZIZSRJK2SnCR24jCoaD/ZpL7yIiT7OnKHCH8PuFE86zRpkx2rCS1yktv1DkvtA
/hE9C7DZVS02t+38WmPvPReepRaLYj0S4PDFP/TxwbrFDOeXnql/PZyyDdfj903m
2FnkdUdlP8B5wVFGijOZp36S9QXRdkC6f/bKdE11XDEyuaw1tJVAQpc+UCHNToX+
28/CKGB4X38FpwxQEcCZhdtcdbcKN+ERGcD+rRmAvxCNov3x/8AuYR3PkmWffGF1
J53Grbmg5rB8Akwz0DjESYg8tpyHxdBKxnY4qHIoSisABtebs0sci90PhAB2w4ua
TaD26tNFDPlqyTDpvpUFvcrcufb7AWkV9HfRxefTKgOkmiSbkAwh+1EZOGwU4OjT
fh8NhVOmfpTycrgF3Ua0/WCXtGOeZAp/9RIyHab0f6C+y59L8TbNRrvMGr/WhWEU
gubigGRGhKrI0FxinGC0n5aoLAb5919ScXTvzQCYnR21j1WC6gSMlkVUZeZVuX2g
SNH7f/liyIEtFlGM8kH0ELtPlhpWorgUrZ5dfSzsECi5J6Dfop31bHwv9JF4p9La
KYN6IrF/LnoOSk4rxTDiEgGPrdNNNvpsJeE8Vx98xvgoAPYoVzgPI2BP5qBbO8wD
ObAAsM6jF1oXr3jhdkUj9ReaMiq7TwrEAmLiAaDyyBzJVzed79I9j9LqZYkkxJhf
0LeaSpCBfSHZ/s3ijQLN9rEEITTgGwJ5YXreiQHcszIFT128AXXPnPOIhcAF2txZ
VWBbxsAHwPyYHhjOaZNCjxuiMFsSEPM4ihsck0FoPqPYoaBqDEHqpdUdywPMFAnj
SWZsNqAdw68IAhIf1H3q1MN96Tr0aF5x1S5H9ZHvr61e8gQxbI0rXG/eRiXVSKwX
3tJwhiYayqjni12FWiUHy2rgZujkbdhtyg3bLvGi3/Qpli8ctaGgOAKgHnLbChDP
Zq+lP4rrlDPQh3p9V/ehtGh0F/7jK5RmeKMjXCsRtonHWL6vZs2G1Eqv4uTVj2eM
ry40k0CLHWUpXMJEP3E1UeDSCYGurHbnqbZrX2SVGdSZNLxkZxuxrfTYRg5ca0tU
Di7IpyqZr7dTGQS3cpnMzUxEdsEyQfQh2uDSUyIlvmlGGY4jDJccHVtKOlg6gBOc
ZTEpzsfhnpakEDPLbWI3xvAssjUkNBbv5+LFA+Z2GeonI7MOyOjAMH2vl4GvoCzA
d8WXjokYaYvEGpmOBrjOJKinz/KNehG3B27EmcaH4laVgRGVd2ivQ+vD/Ydb21r0
92Qxt3jXSDl+cCfT0yJ50cRhH2NhrggDyO3n+EmtGV1GfJUPNMKDznS9S+CNM15U
XwZq0QfhA4qslCgS3vqAVPyNWdLIcc0dIqyr4QtXeiNPSOr8sMKj0H861iYtu5iF
3q7tLg5GAZBvOY9y2uZxtpObZBC1Yz8MD19fy8woLNH8tCaUXRmEOHQ8XtIM3qvd
o34UnFabbKoCSdEpA7/jprnIXp/Qf0iquCFFSCnhrQiAmQj+ETsKRjOwpPQj4NBx
ppwYgvOqpkZsLxGgb+UhR/uoW3r6NkJIFfn2VEc/ofHF3K6cY/sF4ejzCFcEjV5s
eIPmFPVdIhdKzDLLQd1kGsx103SbJwjpfxSB3CFM1ZBdBg2DCuhnQ28Xqbd0HBc1
KXQFDFi4F2+0tUXAbiG7+h2PlXUnC52bMRWE3xE3fXQpgVEmOjB4S6m7QglWSBPL
xp7TSFpFBvCzd2D0L2b+74oS7qppqSc7W0FPHK+Ml5MmoRLhDvp+5jiqqZI4t2Hm
RbJqCz6t3lY9d0+OHRryzqbbZ48wJrDjFzt84Y/s9zAY8QsrkVwegInHTqXzd/mU
moWqN5UuA45gzkAUEy7yFgcOEE8S2XCJkcGtbZtJhFd3EnZE5pvdWEwHUBSbvFrI
zkWw8NvX2QpcGPelim3EMbzncEP/ix/e7/9wvGMQDQlRPsRC4TlsibLRzgfC7B3s
5S4l6S3oIqsz+BM+e6iKONxKjB2BBBfAGvXQ1OXgXv0TE03e3xK+nyt20iZbG7JV
SDwS+VsTXAQ/t8tO+poXpMHyNAQUeYSUxHPJojTWBRH6EzO5whf4vbAH9BuMRaCY
il3KjkeXtU2svZ1nyRD8uNcztLu6b8P7nOGj0+hm1iYDRuwyosJUicLchcumsQjH
SYd35mtF2Mjyje7SXgS06C2uKdNa46cp3sc4I+pc2UETugJnNf2fgckp8liW4PJI
3Pw386i3wCfDyAhRpxD5C+IIITxgPRZ4/D+UnKoh4zB01S7f3lws5x3FFQGL4kmy
iduNHNIaCOgmSd3S5NLOk7natCBZNsSsPjRh3yTutqwblTLYmlFqFF8uWCx9+ae+
T6JT8zJ0Oglz9cqLfEAiHaPCQXsdcPjR2Cf6gAXhaFVvB+Itq/cKEDHtsFfCM6xw
0WM1YeeDIUqcArgr50PuYuuLYBLyKxMqpEDz9F4Bmix1UvYm0ZxD/X94Cyvwq9um
WazkT/OYeFvkPraRxvvXgCCmob275K8fJal8SF1+73cC+rp8DYq99G4urqTW9Rt9
NE25B1gnNsCll+ptRVljVpQmBbo4Wq0kTUgP9eYUapfXje/PGuGE95fNeYoQkQYT
YWrgo/QSdqNB0tSc91CpUY5dDNP4TB/1wWp9lsKAqTwoDbPO3p2fJtPcYSLEX8iw
7V66jYu9+sYYQRgMoT/8DQzJGVU8odOCJ4MespfmM5XYOuGzU/wzwC02MxEwqFix
sx4WDAi9oFo3j9rSa3PSB3IrTUSUAvJMTDrlpWKW1dcPINMXpwYZOyPlvcunPIpS
JIAnfpeb+H58iswhb1r+y4/o7rN4HeV/kautfY5JFC+a6E16H6B5/G8ob6Buzy7Z
S2tMic3gfcKlXqg5gpkkeJed25/J+dSgFoDqHf6yoQxwNY2J5jNgeGph+23QSkcD
Pbi41F7H06DLfPPcJL1aoPRX1eOYOZZzGok1u6P5BYhxPhpOY1e5cDndtQxpnRyt
+W2nAz1ep8N/88aSEBxRj5A3YncfdYopKuOiyrZiCu+0zfQHrcVupJTGSW+clXe3
VLTvpmh2ekzXfhnPZU6lUWTLrtRI+SlKOy8V5Sugiv34eAUxMJxModI4+PQ4Pfba
EFyvp6fri6DvAAkD794ityFnJxiR0MDE2+7HpVvmEy8UDx0We6YsBfdPK1/+3rZA
2z8ue9tOe/2Om34Qg1D18Lj0XNgovvtEuvVrjvU6TuEUc51NDzHUmp5blUtPOIJz
YKwyCcped4PjieY6d+WBzXfSzN+13VDmbA2Izf2pKAx+avYKAXwaQjMzZeInWgNW
F8gynJQD3IrBLXpXFdpPyqWq9BRhnpUOGslyhcxTzS9mlt4SzgX/c91YfEbguCzo
LlJftYFFOPTmJ3mwXUBmnfyVXlssdeWBDaXMN9+XbiJM7dMEVuDg0a+RX+soBKie
+KKewaIqHqSL3PjR4Ln21E8iYo79x3AJogbbYd6WMl/xzoLR0p8xS+tDTCQ8Wmz9
UT9SlStbSMC3jEzHetKd5ZkpEgdfLvk7cJAra149xNEwLd53lUrM8EypKl9l8xrz
7ZCQkhG+OshZC2S79sXLaYAp4BYif7EXMEdIfrBxJlMnW/OZhxx2BWHI2vtBBGIu
2bLTN4R+vqmyp+q6cgUxwRwDIt4aCjSRB81qqrNflh/jFxiC7ZYCUe6nW4PpTjbs
uqokgOs3VZQ0S6RlOltAAXm50+rJyc+PQeStL3RDcNRdIcH8HhUjddwV3l9wARUM
H9KneLcRJTg5dZbs0GpwYxDdy1DIlLbmey51LXEX2JMwpvzy5hlb/LZB0b80zx0q
QSJ2Rs9LRwkHJ38u1zKpYMVRMpbajgOoTrpVbJ5Ex3uzVGozaEPyajxaImAuqX3z
5eHPmpkXF0DYTSj5O59Q7ANvaN8oaT/IMDx/hATnONJgmKexezW9hMDPCKac2dor
ay2kF7YRmBjNMAI3lZAdbPvcZ+M+IIiyvvKJHkSnKFz3Y+ph5BUTFPyZTzvQ2yp0
xmX3y7aChUtnJl79vJsUu0OMjXL8rAA8G0gCD7kXNDeoDRlgeRAK+7+b8VlbQIpf
EjCpwNrpdV0Jn+6lpfn1Tapv7VUQgZChzVYc+4JNRcF0J5fmLz7CVRVYUGbyuxjh
ccTYUz2YitkrZo8S521AB5qvSrYaQNE/VfLiHSDQNbcZth/4lQdh5fCthwrLF6/B
g6sFEM/fykQ7+yUDThPw1CHsnprTRNh+wiDNQ/x3VTXaMf9yxyT3g58Q/BMREoZ8
JlUQO0u0b4rPTfflfy1nK+1c7gxzwZknjmWZ6CxksU+Kxoz9mSYdaEjAohzc24Ue
4KDK2zOx5ja9RFnBIn6S+rWCeRcgns3aHVRqEkVPZYeCVu5U6OllYeGLQ88ihCTL
CIo1sdWdaT9doKxyF9t966XHOJ4vqQietPHsbgGBR2bLAtUmYhIItjffYma4covO
Q5S9RMjqePdt5+Y3Hd7molVUa4v4Rq2hSkZvrvGzLGZ+Cap4CJ8UqUFYMrSNFXdT
Fonk81php4Gq0Dsy0Uq8tJtJ9QDiIWBTcJMC8maiRduj1yUE+XzfSnUihP5wNjho
Z1ETM1lZa17ulqKiVz8jVjTfgXyX34iXDk4oVeyszfc9+dFxka6z4txDuhScOoW7
O6XyF+KBEyXm+/NoeY1Tvn8Hc77pUoXq3Sb7G32RQbXXyizyGgExSnBk5OSi+upq
myDO0+wowmoSx7ENcJ8tZ/I6hxD5Ap5bVZuNi60d+06SjIuES0FPLAB1EkQZI1EB
uY69/+vJv5Mxo2M8IH3uaFY6vbv+kOFxzSKO/TOh97i+2X8GMIy+jld1CZugy/FH
/nDOd6M72LvdxgFL40Ip7WE4BwO5e2ADrgWx5/2TejAf8SbxuyGL7xJ2SqAkiKuw
lPD6yvXKj41kcIGToR9+GWVqtGvoi4FZpNWaUkvtDfcmPe9aSkSiY5oLw2VGcgfM
43zFVUtJhBPK3VaLthn2yl+vVoui9ZUM3XVAsAsC/ZlVOkoiL+of+bysWbRY++3M
iytyRlsxosX+mzErCmJopNVcNE/bUDPKEzSf/ndVAlULbM5TAMitmhvUU8hrL9Fq
HhC2A0RbAdyb58Auxa+/fE9iAUVE/dbx40mmmR9+oWtTx/oAT9tuvO/tErmc3fDz
l2WOoilfq0xdcjvshN5DlZTOR2Qkv0tOzpTbk0JcZ3fyhIMr4dvryphbWsOkICv/
2X6cufjB8IiAbMJyHKWW3VmS7CHs5rwx6sEsO+3Un2j5tI9+1BqmtYZIgQZXmzBV
F6YKSsPCLKm3culSYPGZXd4kBBhdbl8F6UklmoZfpE0pR4vu9oPyjFq6HkZ6lFs9
yXYRcfvPrg6UuTp7rv4oUXlV4sWVzgzH2BnWgCj+nxkHj9HF4LsO7uO7slKJJYjf
bXLDwiHoAtY0SXExYcwkDEV0c3vvh1f1Rtnd2lmqokh7yVMM8VrPgNwhGMRTLXLd
5Ak1V9nTMphrYfPRsUJf8i9uTUBWob2OyU50pT8TiooS6UEj7kIxDOJMSoqYe4IY
SDGfX2vQylsuM60+GYCvWQchFoM6xY/dAw6hA49gwSaeqq5sIMgFAdcsAg+0lits
/B19Mc9WPZVt/KClfducXa2QZmM8lVD+vYlAgZyX1nh0EBhfPX1EG+NRvgPUBp+W
y0aX18uksG65oBqinQBG7+ryGmaLyCcZdJs91nJ+bPpbzG49RoV7uJJ6veua1rqo
ECMFkTtsC9AQ6bIoztBQ97ayYxOcEYSYA7fbF07M/wm+Y24twn/1RU5PGwwwEBwu
5Bha88hIooWfhBy7Mymf9cEbuLeg1yrbs9ImEGdJhZ2V9IebaLB65BR3x6xBUQe2
fgXI+m+uA4lm5My1HVxnFq/ZR/l3+c7yrFDmfyOWdtEm0G4hMh7pdBYx5jp7eUi3
eQVXKM3xWmYgNlR1MLGwVIR3WdaHLm9KTuYW8wBDlCs=
`pragma protect end_protected

//pragma protect end
